module gray_to_bin (
	gray, 
	bin);
   input [6:0] gray;
   output [6:0] bin;

   // Internal wires
   wire FE_PHN682_bin_dout_4_;

   DLY4X1 FE_PHC682_bin_dout_4_ (.Y(bin[4]), 
	.A(FE_PHN682_bin_dout_4_));
   XOR2X1 U1 (.Y(bin[1]), 
	.B(gray[1]), 
	.A(bin[2]));
   XOR2X1 U2 (.Y(bin[5]), 
	.B(gray[6]), 
	.A(gray[5]));
   XOR2X1 U3 (.Y(bin[3]), 
	.B(gray[3]), 
	.A(bin[4]));
   XOR2X1 U4 (.Y(bin[2]), 
	.B(gray[2]), 
	.A(bin[3]));
   XOR2X1 U5 (.Y(FE_PHN682_bin_dout_4_), 
	.B(gray[4]), 
	.A(bin[5]));
   XOR2X1 U6 (.Y(bin[0]), 
	.B(bin[1]), 
	.A(gray[0]));
   BUFX3 U7 (.Y(bin[6]), 
	.A(gray[6]));
endmodule

module control_DW01_inc_0 (
	A, 
	SUM);
   input [6:0] A;
   output [6:0] SUM;

   // Internal wires
   wire FE_PHN3183_bin_dout_6_;
   wire FE_PHN2844_bin_dout_1_;
   wire [6:2] carry;

   BUFXL FE_PHC3183_bin_dout_6_ (.Y(FE_PHN3183_bin_dout_6_), 
	.A(A[6]));
   BUFXL FE_PHC2844_bin_dout_1_ (.Y(FE_PHN2844_bin_dout_1_), 
	.A(A[1]));
   ADDHXL U1_1_5 (.S(SUM[5]), 
	.CO(carry[6]), 
	.B(carry[5]), 
	.A(A[5]));
   ADDHXL U1_1_4 (.S(SUM[4]), 
	.CO(carry[5]), 
	.B(carry[4]), 
	.A(A[4]));
   ADDHXL U1_1_3 (.S(SUM[3]), 
	.CO(carry[4]), 
	.B(carry[3]), 
	.A(A[3]));
   ADDHXL U1_1_2 (.S(SUM[2]), 
	.CO(carry[3]), 
	.B(carry[2]), 
	.A(A[2]));
   ADDHXL U1_1_1 (.S(SUM[1]), 
	.CO(carry[2]), 
	.B(A[0]), 
	.A(FE_PHN2844_bin_dout_1_));
   XOR2X1 U1 (.Y(SUM[6]), 
	.B(FE_PHN3183_bin_dout_6_), 
	.A(carry[6]));
   INVX1 U2 (.Y(SUM[0]), 
	.A(A[0]));
endmodule

module control (
	clk, 
	rst_n, 
	init, 
	next, 
	trig, 
	clk_48Mhz__L6_N43);
   input clk;
   input rst_n;
   output init;
   output next;
   output trig;
   input clk_48Mhz__L6_N43;

   // Internal wires
   wire FE_PHN5059_n21;
   wire FE_PHN2808_init;
   wire FE_PHN822_gray_dout_6_;
   wire FE_PHN753_gray_dout_1_;
   wire FE_PHN752_N7;
   wire FE_PHN681_N8;
   wire FE_PHN678_n20;
   wire FE_PHN536_bin_dout_0_;
   wire FE_PHN534_N9;
   wire FE_PHN439_next;
   wire FE_PHN376_gray_dout_3_;
   wire FE_PHN375_gray_dout_2_;
   wire FE_PHN372_n19;
   wire FE_PHN322_N6;
   wire FE_PHN319_n21;
   wire FE_PHN301_gray_dout_4_;
   wire FE_PHN271_gray_dout_0_;
   wire FE_PHN270_n11;
   wire FE_PHN255_gray_dout_5_;
   wire N4;
   wire N5;
   wire N6;
   wire N7;
   wire N8;
   wire N9;
   wire N10;
   wire n3;
   wire n40;
   wire n50;
   wire n60;
   wire n70;
   wire n80;
   wire n90;
   wire n100;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n1;
   wire n2;
   wire [6:0] bin_dout;
   wire [6:0] bin_add;
   wire [6:0] gray_dout;

   DLY2X1 FE_PHC5059_n21 (.Y(FE_PHN5059_n21), 
	.A(n21));
   DLY2X1 FE_PHC2808_init (.Y(init), 
	.A(FE_PHN2808_init));
   DLY4X1 FE_PHC822_gray_dout_6_ (.Y(FE_PHN822_gray_dout_6_), 
	.A(gray_dout[6]));
   DLY4X1 FE_PHC753_gray_dout_1_ (.Y(FE_PHN753_gray_dout_1_), 
	.A(gray_dout[1]));
   DLY4X1 FE_PHC752_N7 (.Y(FE_PHN752_N7), 
	.A(N7));
   DLY4X1 FE_PHC681_N8 (.Y(FE_PHN681_N8), 
	.A(N8));
   DLY4X1 FE_PHC678_n20 (.Y(FE_PHN678_n20), 
	.A(n20));
   DLY4X1 FE_PHC536_bin_dout_0_ (.Y(FE_PHN536_bin_dout_0_), 
	.A(bin_dout[0]));
   DLY4X1 FE_PHC534_N9 (.Y(FE_PHN534_N9), 
	.A(N9));
   DLY4X1 FE_PHC439_next (.Y(next), 
	.A(FE_PHN439_next));
   DLY4X1 FE_PHC376_gray_dout_3_ (.Y(FE_PHN376_gray_dout_3_), 
	.A(gray_dout[3]));
   DLY4X1 FE_PHC375_gray_dout_2_ (.Y(FE_PHN375_gray_dout_2_), 
	.A(gray_dout[2]));
   DLY4X1 FE_PHC372_n19 (.Y(FE_PHN372_n19), 
	.A(n19));
   DLY4X1 FE_PHC322_N6 (.Y(FE_PHN322_N6), 
	.A(N6));
   DLY4X1 FE_PHC319_n21 (.Y(FE_PHN319_n21), 
	.A(FE_PHN5059_n21));
   DLY4X1 FE_PHC301_gray_dout_4_ (.Y(FE_PHN301_gray_dout_4_), 
	.A(gray_dout[4]));
   DLY4X1 FE_PHC271_gray_dout_0_ (.Y(FE_PHN271_gray_dout_0_), 
	.A(gray_dout[0]));
   DLY4X1 FE_PHC270_n11 (.Y(FE_PHN270_n11), 
	.A(n11));
   DLY4X1 FE_PHC255_gray_dout_5_ (.Y(FE_PHN255_gray_dout_5_), 
	.A(gray_dout[5]));
   DFFRHQX1 next_reg (.RN(rst_n), 
	.Q(FE_PHN439_next), 
	.D(FE_PHN372_n19), 
	.CK(clk));
   DFFRHQX1 gray_dout_reg_0_ (.RN(rst_n), 
	.Q(gray_dout[0]), 
	.D(N4), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 gray_dout_reg_1_ (.RN(rst_n), 
	.Q(gray_dout[1]), 
	.D(N5), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 gray_dout_reg_2_ (.RN(rst_n), 
	.Q(gray_dout[2]), 
	.D(FE_PHN322_N6), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 gray_dout_reg_5_ (.RN(rst_n), 
	.Q(gray_dout[5]), 
	.D(FE_PHN534_N9), 
	.CK(clk));
   DFFRHQX1 gray_dout_reg_4_ (.RN(rst_n), 
	.Q(gray_dout[4]), 
	.D(FE_PHN681_N8), 
	.CK(clk));
   DFFRHQX1 gray_dout_reg_6_ (.RN(rst_n), 
	.Q(gray_dout[6]), 
	.D(N10), 
	.CK(clk));
   DFFRHQX1 gray_dout_reg_3_ (.RN(rst_n), 
	.Q(gray_dout[3]), 
	.D(FE_PHN752_N7), 
	.CK(clk));
   DFFRHQX1 init_reg (.RN(rst_n), 
	.Q(FE_PHN2808_init), 
	.D(FE_PHN678_n20), 
	.CK(clk));
   DFFRHQX1 trig_reg (.RN(rst_n), 
	.Q(trig), 
	.D(FE_PHN319_n21), 
	.CK(clk));
   NOR2X1 U3 (.Y(N9), 
	.B(n12), 
	.A(FE_PHN270_n11));
   XNOR2X1 U4 (.Y(n12), 
	.B(bin_add[6]), 
	.A(bin_add[5]));
   NOR2X1 U5 (.Y(N8), 
	.B(n13), 
	.A(FE_PHN270_n11));
   XNOR2X1 U6 (.Y(n13), 
	.B(bin_add[5]), 
	.A(bin_add[4]));
   NOR2BX1 U7 (.Y(N10), 
	.B(FE_PHN270_n11), 
	.AN(bin_add[6]));
   NOR2X1 U8 (.Y(N7), 
	.B(n14), 
	.A(FE_PHN270_n11));
   XNOR2X1 U9 (.Y(n14), 
	.B(bin_add[4]), 
	.A(bin_add[3]));
   NOR2X1 U10 (.Y(N6), 
	.B(n15), 
	.A(FE_PHN270_n11));
   XNOR2X1 U11 (.Y(n15), 
	.B(bin_add[3]), 
	.A(bin_add[2]));
   NOR2X1 U12 (.Y(N5), 
	.B(n16), 
	.A(FE_PHN270_n11));
   XNOR2X1 U13 (.Y(n16), 
	.B(bin_add[2]), 
	.A(bin_add[1]));
   NOR2X1 U14 (.Y(N4), 
	.B(n17), 
	.A(FE_PHN270_n11));
   XNOR2X1 U15 (.Y(n17), 
	.B(bin_add[0]), 
	.A(bin_add[1]));
   NAND3X1 U16 (.Y(n3), 
	.C(FE_PHN375_gray_dout_2_), 
	.B(FE_PHN376_gray_dout_3_), 
	.A(FE_PHN271_gray_dout_0_));
   INVX1 U17 (.Y(n1), 
	.A(FE_PHN271_gray_dout_0_));
   OAI2BB2X1 U18 (.Y(n19), 
	.B1(n40), 
	.B0(n3), 
	.A1N(n40), 
	.A0N(next));
   NAND4X1 U19 (.Y(n40), 
	.D(n60), 
	.C(n50), 
	.B(FE_PHN375_gray_dout_2_), 
	.A(FE_PHN301_gray_dout_4_));
   NOR3X1 U20 (.Y(n60), 
	.C(FE_PHN255_gray_dout_5_), 
	.B(FE_PHN822_gray_dout_6_), 
	.A(FE_PHN753_gray_dout_1_));
   XNOR2X1 U21 (.Y(n50), 
	.B(FE_PHN376_gray_dout_3_), 
	.A(FE_PHN271_gray_dout_0_));
   OAI2BB2X1 U22 (.Y(n20), 
	.B1(n70), 
	.B0(n3), 
	.A1N(n70), 
	.A0N(init));
   NAND3X1 U23 (.Y(n70), 
	.C(n80), 
	.B(FE_PHN376_gray_dout_3_), 
	.A(FE_PHN375_gray_dout_2_));
   OAI2BB2X1 U24 (.Y(n21), 
	.B1(n90), 
	.B0(n1), 
	.A1N(n90), 
	.A0N(trig));
   NAND3BX1 U25 (.Y(n90), 
	.C(n80), 
	.B(n2), 
	.AN(FE_PHN375_gray_dout_2_));
   INVX1 U26 (.Y(n2), 
	.A(FE_PHN376_gray_dout_3_));
   AND4X2 U27 (.Y(n11), 
	.D(FE_PHN753_gray_dout_1_), 
	.C(n18), 
	.B(FE_PHN255_gray_dout_5_), 
	.A(FE_PHN822_gray_dout_6_));
   NOR2BX1 U28 (.Y(n18), 
	.B(n3), 
	.AN(FE_PHN301_gray_dout_4_));
   NOR4BX1 U29 (.Y(n80), 
	.D(FE_PHN822_gray_dout_6_), 
	.C(FE_PHN255_gray_dout_5_), 
	.B(FE_PHN301_gray_dout_4_), 
	.AN(n100));
   XNOR2X1 U30 (.Y(n100), 
	.B(n1), 
	.A(FE_PHN753_gray_dout_1_));
   gray_to_bin gtb (.gray({ FE_PHN822_gray_dout_6_,
		FE_PHN255_gray_dout_5_,
		FE_PHN301_gray_dout_4_,
		FE_PHN376_gray_dout_3_,
		FE_PHN375_gray_dout_2_,
		FE_PHN753_gray_dout_1_,
		FE_PHN271_gray_dout_0_ }), 
	.bin(bin_dout));
   control_DW01_inc_0 add_15 (.A({ bin_dout[6],
		bin_dout[5],
		bin_dout[4],
		bin_dout[3],
		bin_dout[2],
		bin_dout[1],
		FE_PHN536_bin_dout_0_ }), 
	.SUM(bin_add));
endmodule

module aes_encipher_block (
	clk, 
	reset_n, 
	next, 
	round, 
	round_key, 
	sboxw, 
	new_sboxw, 
	block, 
	new_block, 
	ready, 
	FE_OFN39_reset_n, 
	FE_OFN43_reset_n, 
	FE_OFN49_reset_n, 
	FE_OFN50_reset_n, 
	FE_OFN51_reset_n, 
	FE_OFN54_reset_n, 
	FE_OFN55_reset_n, 
	FE_OFN56_reset_n, 
	clk_48Mhz__L6_N23, 
	clk_48Mhz__L6_N37, 
	clk_48Mhz__L6_N39, 
	clk_48Mhz__L6_N40, 
	clk_48Mhz__L6_N41, 
	clk_48Mhz__L6_N44, 
	clk_48Mhz__L6_N46, 
	clk_48Mhz__L6_N47, 
	clk_48Mhz__L6_N5, 
	clk_48Mhz__L6_N8, 
	clk_48Mhz__L6_N9);
   input clk;
   input reset_n;
   input next;
   output [3:0] round;
   input [127:0] round_key;
   output [31:0] sboxw;
   input [31:0] new_sboxw;
   input [127:0] block;
   output [127:0] new_block;
   output ready;
   input FE_OFN39_reset_n;
   input FE_OFN43_reset_n;
   input FE_OFN49_reset_n;
   input FE_OFN50_reset_n;
   input FE_OFN51_reset_n;
   input FE_OFN54_reset_n;
   input FE_OFN55_reset_n;
   input FE_OFN56_reset_n;
   input clk_48Mhz__L6_N23;
   input clk_48Mhz__L6_N37;
   input clk_48Mhz__L6_N39;
   input clk_48Mhz__L6_N40;
   input clk_48Mhz__L6_N41;
   input clk_48Mhz__L6_N44;
   input clk_48Mhz__L6_N46;
   input clk_48Mhz__L6_N47;
   input clk_48Mhz__L6_N5;
   input clk_48Mhz__L6_N8;
   input clk_48Mhz__L6_N9;

   // Internal wires
   wire FE_PHN5256_n892;
   wire FE_PHN5253_n1256;
   wire FE_PHN5252_n1296;
   wire FE_PHN5251_n866;
   wire FE_PHN5250_n1264;
   wire FE_PHN5249_n1331;
   wire FE_PHN5248_n1236;
   wire FE_PHN5247_n1268;
   wire FE_PHN5246_n1276;
   wire FE_PHN5245_n1240;
   wire FE_PHN5244_n1138;
   wire FE_PHN5235_n658;
   wire FE_PHN5233_n929;
   wire FE_PHN5229_n1274;
   wire FE_PHN5228_n782;
   wire FE_PHN5227_n1256;
   wire FE_PHN5226_n1241;
   wire FE_PHN5225_n1238;
   wire FE_PHN5224_n541;
   wire FE_PHN5223_n1292;
   wire FE_PHN5222_n1283;
   wire FE_PHN5221_n323;
   wire FE_PHN5220_n1227;
   wire FE_PHN5219_n1252;
   wire FE_PHN5218_n1279;
   wire FE_PHN5217_n1266;
   wire FE_PHN5216_n1244;
   wire FE_PHN5215_n1329;
   wire FE_PHN5214_n774;
   wire FE_PHN5213_n1138;
   wire FE_PHN5212_n1296;
   wire FE_PHN5211_n1331;
   wire FE_PHN5210_n1264;
   wire FE_PHN5209_n1236;
   wire FE_PHN5208_n1240;
   wire FE_PHN5207_n866;
   wire FE_PHN5206_n316;
   wire FE_PHN5205_n1273;
   wire FE_PHN5204_n1229;
   wire FE_PHN5203_n1209;
   wire FE_PHN5202_n1272;
   wire FE_PHN5201_n1225;
   wire FE_PHN5200_n1249;
   wire FE_PHN5199_n1268;
   wire FE_PHN5198_n1208;
   wire FE_PHN5197_n1276;
   wire FE_PHN5196_n1270;
   wire FE_PHN5195_n1289;
   wire FE_PHN5194_n1328;
   wire FE_PHN5193_n1291;
   wire FE_PHN5192_n1265;
   wire FE_PHN5191_n1257;
   wire FE_PHN5190_n1280;
   wire FE_PHN5189_n1248;
   wire FE_PHN5188_n1218;
   wire FE_PHN5187_n1233;
   wire FE_PHN5186_n1247;
   wire FE_PHN5185_n1235;
   wire FE_PHN5184_n1219;
   wire FE_PHN5183_n1282;
   wire FE_PHN5182_n1242;
   wire FE_PHN5181_n1326;
   wire FE_PHN5180_n1297;
   wire FE_PHN5179_n1269;
   wire FE_PHN5178_n1239;
   wire FE_PHN5177_n1324;
   wire FE_PHN5176_n1234;
   wire FE_PHN5175_n1250;
   wire FE_PHN5174_n1232;
   wire FE_PHN5172_n1100;
   wire FE_PHN5169_n1297;
   wire FE_PHN5168_n1072;
   wire FE_PHN5167_n1028;
   wire FE_PHN5166_n1219;
   wire FE_PHN5165_n563;
   wire FE_PHN5164_n1131;
   wire FE_PHN5163_n1291;
   wire FE_PHN5162_n1274;
   wire FE_PHN5161_n426;
   wire FE_PHN5160_n1307;
   wire FE_PHN5153_n1265;
   wire FE_PHN5152_n1090;
   wire FE_PHN5151_n1283;
   wire FE_PHN5150_n782;
   wire FE_PHN5149_n1240;
   wire FE_PHN5148_n372;
   wire FE_PHN5147_n1219;
   wire FE_PHN5146_n548;
   wire FE_PHN5145_n1302;
   wire FE_PHN5144_n1078;
   wire FE_PHN5143_n1305;
   wire FE_PHN5142_n309;
   wire FE_PHN5141_n1257;
   wire FE_PHN5140_n1206;
   wire FE_PHN5139_n1239;
   wire FE_PHN5138_n1250;
   wire FE_PHN5137_n1072;
   wire FE_PHN5136_n1251;
   wire FE_PHN5135_n1237;
   wire FE_PHN5134_n541;
   wire FE_PHN5133_n1043;
   wire FE_PHN5132_n378;
   wire FE_PHN5131_n1300;
   wire FE_PHN5130_n1210;
   wire FE_PHN5129_n1307;
   wire FE_PHN5128_n426;
   wire FE_PHN5127_n1035;
   wire FE_PHN5126_n1021;
   wire FE_PHN5125_n366;
   wire FE_PHN5124_n1212;
   wire FE_PHN5123_n1323;
   wire FE_PHN5122_n1213;
   wire FE_PHN5121_n1314;
   wire FE_PHN5120_n1230;
   wire FE_PHN5119_n651;
   wire FE_PHN5118_n1308;
   wire FE_PHN5117_n1274;
   wire FE_PHN5116_n1322;
   wire FE_PHN5115_n1303;
   wire FE_PHN5114_n1276;
   wire FE_PHN5113_n1242;
   wire FE_PHN5112_n1028;
   wire FE_PHN5111_n1275;
   wire FE_PHN5110_n441;
   wire FE_PHN5109_n696;
   wire FE_PHN5108_n1241;
   wire FE_PHN5107_n1220;
   wire FE_PHN5106_n1315;
   wire FE_PHN5105_n1269;
   wire FE_PHN5104_n1297;
   wire FE_PHN5103_n563;
   wire FE_PHN5102_n1131;
   wire FE_PHN5101_n1066;
   wire FE_PHN5100_n1244;
   wire FE_PHN5099_n1243;
   wire FE_PHN5098_n1282;
   wire FE_PHN5097_n1333;
   wire FE_PHN5096_n1221;
   wire FE_PHN5095_n1211;
   wire FE_PHN5094_n1267;
   wire FE_PHN5093_n1236;
   wire FE_PHN5092_n1291;
   wire FE_PHN5091_n1098;
   wire FE_PHN5090_n1306;
   wire FE_PHN5089_n1324;
   wire FE_PHN5088_n1281;
   wire FE_PHN5087_n1304;
   wire FE_PHN5086_n1266;
   wire FE_PHN5085_n1233;
   wire FE_PHN5084_n1226;
   wire FE_PHN5083_n1228;
   wire FE_PHN5082_n1245;
   wire FE_PHN5081_n1290;
   wire FE_PHN5080_n1235;
   wire FE_PHN5079_n1299;
   wire FE_PHN5078_n1258;
   wire FE_PHN5075_n419;
   wire FE_PHN5045_n1334;
   wire FE_PHN3408_enc_ctrl_reg_0_;
   wire FE_PHN3108_Dout_104_;
   wire FE_PHN3107_Dout_33_;
   wire FE_PHN3106_Dout_97_;
   wire FE_PHN3105_Dout_47_;
   wire FE_PHN3104_Dout_8_;
   wire FE_PHN3095_Dout_119_;
   wire FE_PHN3081_n1194;
   wire FE_PHN2856_n1338;
   wire FE_PHN2850_Dout_125_;
   wire FE_PHN2843_n1335;
   wire FE_PHN2821_enc_ctrl_reg_1_;
   wire FE_PHN2816_n1013;
   wire FE_PHN2813_enc_round_nr_2_;
   wire FE_PHN2812_enc_round_nr_1_;
   wire FE_PHN2809_n1340;
   wire FE_PHN2807_n1330;
   wire FE_PHN2806_n1301;
   wire FE_PHN2805_n1227;
   wire FE_PHN1310_n1334;
   wire FE_PHN821_Dout_1_;
   wire FE_PHN751_n1337;
   wire FE_PHN750_Dout_103_;
   wire FE_PHN703_n1336;
   wire FE_PHN702_Dout_38_;
   wire FE_PHN701_Dout_36_;
   wire FE_PHN604_Dout_34_;
   wire FE_PHN603_Dout_10_;
   wire FE_PHN602_n1197;
   wire FE_PHN601_Dout_46_;
   wire FE_PHN600_Dout_37_;
   wire FE_PHN599_Dout_102_;
   wire FE_PHN598_Dout_116_;
   wire FE_PHN597_Dout_44_;
   wire FE_PHN596_Dout_101_;
   wire FE_PHN595_Dout_110_;
   wire FE_PHN535_enc_ctrl_we;
   wire FE_PHN533_Dout_122_;
   wire FE_PHN528_Dout_111_;
   wire FE_PHN444_Dout_73_;
   wire FE_PHN443_Dout_72_;
   wire FE_PHN442_Dout_114_;
   wire FE_PHN441_Dout_9_;
   wire FE_PHN440_Dout_54_;
   wire FE_PHN438_Dout_0_;
   wire FE_PHN437_Dout_108_;
   wire FE_PHN436_Dout_117_;
   wire FE_PHN435_Dout_109_;
   wire FE_PHN433_Dout_100_;
   wire FE_PHN415_Dout_93_;
   wire FE_PHN414_Dout_63_;
   wire FE_PHN413_Dout_120_;
   wire FE_PHN412_Dout_126_;
   wire FE_PHN410_enc_ctrl_reg_0_;
   wire FE_PHN378_Dout_39_;
   wire FE_PHN377_Dout_6_;
   wire FE_PHN374_Dout_53_;
   wire FE_PHN373_Dout_68_;
   wire FE_PHN371_Dout_35_;
   wire FE_PHN369_Dout_105_;
   wire FE_PHN368_Dout_74_;
   wire FE_PHN367_Dout_76_;
   wire FE_PHN366_Dout_20_;
   wire FE_PHN365_Dout_22_;
   wire FE_PHN364_Dout_21_;
   wire FE_PHN363_Dout_3_;
   wire FE_PHN362_Dout_45_;
   wire FE_PHN361_Dout_127_;
   wire FE_PHN356_Dout_26_;
   wire FE_PHN355_Dout_58_;
   wire FE_PHN354_n1335;
   wire FE_PHN353_Dout_60_;
   wire FE_PHN352_Dout_123_;
   wire FE_PHN351_Dout_121_;
   wire FE_PHN350_Dout_124_;
   wire FE_PHN341_Dout_79_;
   wire FE_PHN340_Dout_65_;
   wire FE_PHN339_Dout_107_;
   wire FE_PHN338_Dout_11_;
   wire FE_PHN337_Dout_115_;
   wire FE_PHN336_Dout_15_;
   wire FE_PHN335_Dout_112_;
   wire FE_PHN334_Dout_49_;
   wire FE_PHN333_Dout_48_;
   wire FE_PHN332_Dout_52_;
   wire FE_PHN331_Dout_17_;
   wire FE_PHN330_Dout_118_;
   wire FE_PHN329_Dout_4_;
   wire FE_PHN328_Dout_113_;
   wire FE_PHN321_Dout_90_;
   wire FE_PHN320_Dout_88_;
   wire FE_PHN318_Dout_62_;
   wire FE_PHN317_Dout_19_;
   wire FE_PHN316_Dout_85_;
   wire FE_PHN315_Dout_42_;
   wire FE_PHN314_Dout_18_;
   wire FE_PHN313_Dout_32_;
   wire FE_PHN312_Dout_50_;
   wire FE_PHN311_Dout_99_;
   wire FE_PHN310_Dout_16_;
   wire FE_PHN309_Dout_70_;
   wire FE_PHN308_Dout_80_;
   wire FE_PHN307_Dout_13_;
   wire FE_PHN306_Dout_51_;
   wire FE_PHN305_Dout_41_;
   wire FE_PHN304_Dout_95_;
   wire FE_PHN303_Dout_92_;
   wire FE_PHN302_Dout_28_;
   wire FE_PHN300_Dout_55_;
   wire FE_PHN299_Dout_23_;
   wire FE_PHN298_Dout_7_;
   wire FE_PHN297_Dout_64_;
   wire FE_PHN296_Dout_84_;
   wire FE_PHN295_Dout_14_;
   wire FE_PHN294_Dout_77_;
   wire FE_PHN293_Dout_75_;
   wire FE_PHN292_Dout_78_;
   wire FE_PHN289_Dout_91_;
   wire FE_PHN288_Dout_94_;
   wire FE_PHN287_Dout_59_;
   wire FE_PHN286_Dout_24_;
   wire FE_PHN285_Dout_25_;
   wire FE_PHN284_Dout_57_;
   wire FE_PHN282_Dout_30_;
   wire FE_PHN281_Dout_31_;
   wire FE_PHN280_Dout_40_;
   wire FE_PHN279_Dout_86_;
   wire FE_PHN278_Dout_87_;
   wire FE_PHN277_Dout_81_;
   wire FE_PHN276_Dout_67_;
   wire FE_PHN275_Dout_12_;
   wire FE_PHN274_Dout_82_;
   wire FE_PHN273_Dout_66_;
   wire FE_PHN272_Dout_89_;
   wire FE_PHN269_Dout_71_;
   wire FE_PHN268_Dout_96_;
   wire FE_PHN267_Dout_83_;
   wire FE_PHN266_Dout_98_;
   wire FE_PHN264_Dout_27_;
   wire FE_PHN263_Dout_56_;
   wire FE_PHN262_Dout_61_;
   wire FE_PHN261_Dout_69_;
   wire FE_PHN260_Dout_43_;
   wire FE_PHN259_Dout_5_;
   wire FE_PHN258_n1339;
   wire FE_PHN257_Dout_29_;
   wire FE_PHN256_n943;
   wire FE_PHN253_n704;
   wire FE_PHN252_n1221;
   wire FE_PHN251_n1229;
   wire FE_PHN250_n1223;
   wire FE_PHN249_n1222;
   wire FE_PHN248_n1316;
   wire FE_PHN247_n1332;
   wire FE_PHN246_n1317;
   wire FE_PHN245_n1324;
   wire FE_PHN244_n1322;
   wire FE_PHN243_n1224;
   wire FE_PHN242_n1318;
   wire FE_PHN241_n1252;
   wire FE_PHN240_n1287;
   wire FE_PHN239_n1284;
   wire FE_PHN238_n1319;
   wire FE_PHN237_n1254;
   wire FE_PHN236_n1292;
   wire FE_PHN235_n1285;
   wire FE_PHN234_n1255;
   wire FE_PHN233_n1253;
   wire FE_PHN232_n1286;
   wire FE_PHN231_n1227;
   wire FE_PHN230_n1290;
   wire FE_PHN229_n1216;
   wire FE_PHN228_n1300;
   wire FE_PHN227_n1258;
   wire FE_PHN226_n1214;
   wire FE_PHN225_n1277;
   wire FE_PHN224_n1327;
   wire FE_PHN223_n1228;
   wire FE_PHN222_n1215;
   wire FE_PHN221_n1309;
   wire FE_PHN220_n1311;
   wire FE_PHN219_n1232;
   wire FE_PHN218_n1226;
   wire FE_PHN217_n1295;
   wire FE_PHN216_n1260;
   wire FE_PHN215_n1323;
   wire FE_PHN214_n1310;
   wire FE_PHN213_n1330;
   wire FE_PHN212_n1246;
   wire FE_PHN211_n1289;
   wire FE_PHN210_n1314;
   wire FE_PHN209_n1250;
   wire FE_PHN208_n1245;
   wire FE_PHN207_n1247;
   wire FE_PHN206_n1333;
   wire FE_PHN205_n1282;
   wire FE_PHN204_n1235;
   wire FE_PHN203_n1291;
   wire FE_PHN202_n1325;
   wire FE_PHN201_n1219;
   wire FE_PHN200_n1298;
   wire FE_PHN199_n1326;
   wire FE_PHN197_n1320;
   wire FE_PHN196_n1279;
   wire FE_PHN195_n1278;
   wire FE_PHN194_n1256;
   wire FE_PHN193_n1263;
   wire FE_PHN192_n1294;
   wire FE_PHN191_n1293;
   wire FE_PHN190_n1242;
   wire FE_PHN189_n1329;
   wire FE_PHN188_n1331;
   wire FE_PHN187_n1313;
   wire FE_PHN186_n1321;
   wire FE_PHN185_n1312;
   wire FE_PHN184_n1217;
   wire FE_PHN183_n1225;
   wire FE_PHN182_n1236;
   wire FE_PHN181_n1266;
   wire FE_PHN180_n1230;
   wire FE_PHN179_n1234;
   wire FE_PHN177_n1220;
   wire FE_PHN176_n1315;
   wire FE_PHN175_n1283;
   wire FE_PHN174_n1251;
   wire FE_PHN173_n1249;
   wire FE_PHN172_n1218;
   wire FE_PHN171_n1288;
   wire FE_PHN170_n1262;
   wire FE_PHN169_n1248;
   wire FE_PHN168_n1261;
   wire FE_PHN167_n1299;
   wire FE_PHN166_n1328;
   wire FE_PHN165_n1281;
   wire FE_PHN164_n1233;
   wire FE_PHN163_n1280;
   wire FE_PHN162_n1244;
   wire FE_PHN161_n1297;
   wire FE_PHN160_n1267;
   wire FE_PHN159_n1265;
   wire FE_PHN158_n1264;
   wire FE_PHN157_n237;
   wire FE_PHN156_n1213;
   wire FE_PHN154_n1308;
   wire FE_PHN153_n1276;
   wire FE_PHN152_n1237;
   wire FE_PHN151_n1296;
   wire FE_PHN150_n1257;
   wire FE_PHN149_n1259;
   wire FE_PHN148_n1239;
   wire FE_PHN147_n1207;
   wire FE_PHN146_n1206;
   wire FE_PHN145_n1238;
   wire FE_PHN144_n1269;
   wire FE_PHN143_n1302;
   wire FE_PHN142_n1304;
   wire FE_PHN141_n1301;
   wire FE_PHN140_n1208;
   wire FE_PHN139_n1303;
   wire FE_PHN138_n1270;
   wire FE_PHN137_n1271;
   wire FE_PHN136_n1231;
   wire FE_PHN135_n1274;
   wire FE_PHN134_n1211;
   wire FE_PHN133_n1241;
   wire FE_PHN132_n1243;
   wire FE_PHN131_n1240;
   wire FE_PHN130_n1209;
   wire FE_PHN129_n1192;
   wire FE_PHN128_n1275;
   wire FE_PHN127_n1307;
   wire FE_PHN126_n1210;
   wire FE_PHN125_n1305;
   wire FE_PHN123_n1273;
   wire FE_PHN122_n1306;
   wire FE_PHN121_n1212;
   wire FE_PHN118_n1272;
   wire FE_PHN117_n1268;
   wire FE_PHN114_sword_ctr_reg_1_;
   wire FE_PHN113_n1189;
   wire FE_PHN111_enc_ctrl_reg_1_;
   wire FE_OFN98_n232;
   wire FE_OFN97_n232;
   wire enc_ctrl_we;
   wire n54;
   wire n56;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire n478;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire n556;
   wire n557;
   wire n558;
   wire n559;
   wire n560;
   wire n561;
   wire n562;
   wire n563;
   wire n564;
   wire n565;
   wire n566;
   wire n567;
   wire n568;
   wire n569;
   wire n570;
   wire n571;
   wire n572;
   wire n573;
   wire n574;
   wire n575;
   wire n576;
   wire n577;
   wire n578;
   wire n579;
   wire n580;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire n593;
   wire n594;
   wire n595;
   wire n596;
   wire n597;
   wire n598;
   wire n599;
   wire n600;
   wire n601;
   wire n602;
   wire n603;
   wire n604;
   wire n605;
   wire n606;
   wire n607;
   wire n608;
   wire n609;
   wire n610;
   wire n611;
   wire n612;
   wire n613;
   wire n614;
   wire n615;
   wire n616;
   wire n617;
   wire n618;
   wire n619;
   wire n620;
   wire n621;
   wire n622;
   wire n623;
   wire n624;
   wire n625;
   wire n626;
   wire n627;
   wire n628;
   wire n629;
   wire n630;
   wire n631;
   wire n632;
   wire n633;
   wire n634;
   wire n635;
   wire n636;
   wire n637;
   wire n638;
   wire n639;
   wire n640;
   wire n641;
   wire n642;
   wire n643;
   wire n644;
   wire n645;
   wire n646;
   wire n647;
   wire n648;
   wire n649;
   wire n650;
   wire n651;
   wire n652;
   wire n653;
   wire n654;
   wire n655;
   wire n656;
   wire n657;
   wire n658;
   wire n659;
   wire n660;
   wire n661;
   wire n662;
   wire n663;
   wire n664;
   wire n665;
   wire n666;
   wire n667;
   wire n668;
   wire n669;
   wire n670;
   wire n671;
   wire n672;
   wire n673;
   wire n674;
   wire n675;
   wire n676;
   wire n677;
   wire n678;
   wire n679;
   wire n680;
   wire n681;
   wire n682;
   wire n683;
   wire n684;
   wire n685;
   wire n686;
   wire n687;
   wire n688;
   wire n689;
   wire n690;
   wire n691;
   wire n692;
   wire n693;
   wire n694;
   wire n695;
   wire n696;
   wire n697;
   wire n698;
   wire n699;
   wire n700;
   wire n701;
   wire n702;
   wire n703;
   wire n704;
   wire n706;
   wire n707;
   wire n708;
   wire n709;
   wire n710;
   wire n711;
   wire n712;
   wire n713;
   wire n714;
   wire n715;
   wire n716;
   wire n717;
   wire n718;
   wire n719;
   wire n720;
   wire n721;
   wire n722;
   wire n723;
   wire n724;
   wire n725;
   wire n726;
   wire n727;
   wire n728;
   wire n729;
   wire n730;
   wire n731;
   wire n732;
   wire n733;
   wire n734;
   wire n735;
   wire n736;
   wire n737;
   wire n738;
   wire n739;
   wire n740;
   wire n741;
   wire n742;
   wire n743;
   wire n744;
   wire n745;
   wire n746;
   wire n747;
   wire n748;
   wire n749;
   wire n750;
   wire n751;
   wire n752;
   wire n753;
   wire n754;
   wire n755;
   wire n756;
   wire n757;
   wire n758;
   wire n759;
   wire n760;
   wire n761;
   wire n762;
   wire n763;
   wire n764;
   wire n765;
   wire n766;
   wire n767;
   wire n768;
   wire n769;
   wire n770;
   wire n771;
   wire n772;
   wire n773;
   wire n774;
   wire n775;
   wire n776;
   wire n777;
   wire n778;
   wire n779;
   wire n780;
   wire n781;
   wire n782;
   wire n783;
   wire n784;
   wire n785;
   wire n786;
   wire n787;
   wire n788;
   wire n789;
   wire n790;
   wire n791;
   wire n792;
   wire n793;
   wire n794;
   wire n795;
   wire n796;
   wire n797;
   wire n798;
   wire n799;
   wire n800;
   wire n801;
   wire n802;
   wire n803;
   wire n804;
   wire n805;
   wire n806;
   wire n807;
   wire n808;
   wire n809;
   wire n810;
   wire n811;
   wire n812;
   wire n813;
   wire n814;
   wire n815;
   wire n816;
   wire n817;
   wire n818;
   wire n819;
   wire n820;
   wire n821;
   wire n822;
   wire n823;
   wire n824;
   wire n825;
   wire n826;
   wire n827;
   wire n828;
   wire n829;
   wire n830;
   wire n831;
   wire n832;
   wire n833;
   wire n834;
   wire n835;
   wire n836;
   wire n837;
   wire n838;
   wire n839;
   wire n840;
   wire n841;
   wire n842;
   wire n843;
   wire n844;
   wire n845;
   wire n846;
   wire n847;
   wire n848;
   wire n849;
   wire n850;
   wire n851;
   wire n852;
   wire n853;
   wire n854;
   wire n855;
   wire n856;
   wire n857;
   wire n858;
   wire n859;
   wire n860;
   wire n861;
   wire n862;
   wire n863;
   wire n864;
   wire n865;
   wire n866;
   wire n867;
   wire n868;
   wire n869;
   wire n870;
   wire n871;
   wire n872;
   wire n873;
   wire n874;
   wire n875;
   wire n876;
   wire n877;
   wire n878;
   wire n879;
   wire n880;
   wire n881;
   wire n882;
   wire n883;
   wire n884;
   wire n885;
   wire n886;
   wire n887;
   wire n888;
   wire n889;
   wire n890;
   wire n891;
   wire n892;
   wire n893;
   wire n894;
   wire n895;
   wire n896;
   wire n897;
   wire n898;
   wire n899;
   wire n900;
   wire n901;
   wire n902;
   wire n903;
   wire n904;
   wire n905;
   wire n906;
   wire n907;
   wire n908;
   wire n909;
   wire n910;
   wire n911;
   wire n912;
   wire n913;
   wire n914;
   wire n915;
   wire n916;
   wire n917;
   wire n918;
   wire n919;
   wire n920;
   wire n921;
   wire n922;
   wire n923;
   wire n924;
   wire n925;
   wire n926;
   wire n927;
   wire n928;
   wire n929;
   wire n930;
   wire n931;
   wire n932;
   wire n933;
   wire n934;
   wire n935;
   wire n936;
   wire n937;
   wire n938;
   wire n939;
   wire n940;
   wire n941;
   wire n942;
   wire n943;
   wire n945;
   wire n946;
   wire n947;
   wire n948;
   wire n949;
   wire n950;
   wire n951;
   wire n952;
   wire n953;
   wire n954;
   wire n955;
   wire n956;
   wire n957;
   wire n958;
   wire n959;
   wire n960;
   wire n961;
   wire n962;
   wire n963;
   wire n964;
   wire n965;
   wire n966;
   wire n967;
   wire n968;
   wire n969;
   wire n970;
   wire n971;
   wire n972;
   wire n973;
   wire n974;
   wire n975;
   wire n976;
   wire n977;
   wire n978;
   wire n979;
   wire n980;
   wire n981;
   wire n982;
   wire n983;
   wire n984;
   wire n985;
   wire n986;
   wire n987;
   wire n988;
   wire n989;
   wire n990;
   wire n991;
   wire n992;
   wire n993;
   wire n994;
   wire n995;
   wire n996;
   wire n997;
   wire n998;
   wire n999;
   wire n1000;
   wire n1001;
   wire n1002;
   wire n1003;
   wire n1004;
   wire n1005;
   wire n1006;
   wire n1007;
   wire n1008;
   wire n1009;
   wire n1010;
   wire n1011;
   wire n1012;
   wire n1013;
   wire n1014;
   wire n1015;
   wire n1016;
   wire n1017;
   wire n1018;
   wire n1019;
   wire n1020;
   wire n1021;
   wire n1022;
   wire n1023;
   wire n1024;
   wire n1025;
   wire n1026;
   wire n1027;
   wire n1028;
   wire n1029;
   wire n1030;
   wire n1031;
   wire n1032;
   wire n1033;
   wire n1034;
   wire n1035;
   wire n1036;
   wire n1037;
   wire n1038;
   wire n1039;
   wire n1040;
   wire n1041;
   wire n1042;
   wire n1043;
   wire n1044;
   wire n1045;
   wire n1046;
   wire n1047;
   wire n1048;
   wire n1049;
   wire n1050;
   wire n1051;
   wire n1052;
   wire n1053;
   wire n1054;
   wire n1055;
   wire n1056;
   wire n1057;
   wire n1058;
   wire n1059;
   wire n1060;
   wire n1061;
   wire n1062;
   wire n1063;
   wire n1064;
   wire n1065;
   wire n1066;
   wire n1067;
   wire n1068;
   wire n1069;
   wire n1070;
   wire n1071;
   wire n1072;
   wire n1073;
   wire n1074;
   wire n1075;
   wire n1076;
   wire n1077;
   wire n1078;
   wire n1079;
   wire n1080;
   wire n1081;
   wire n1082;
   wire n1083;
   wire n1084;
   wire n1085;
   wire n1086;
   wire n1087;
   wire n1088;
   wire n1089;
   wire n1090;
   wire n1091;
   wire n1092;
   wire n1093;
   wire n1094;
   wire n1095;
   wire n1096;
   wire n1097;
   wire n1098;
   wire n1099;
   wire n1100;
   wire n1101;
   wire n1102;
   wire n1103;
   wire n1104;
   wire n1105;
   wire n1106;
   wire n1107;
   wire n1108;
   wire n1109;
   wire n1110;
   wire n1111;
   wire n1112;
   wire n1113;
   wire n1114;
   wire n1115;
   wire n1116;
   wire n1117;
   wire n1118;
   wire n1119;
   wire n1120;
   wire n1121;
   wire n1122;
   wire n1123;
   wire n1124;
   wire n1125;
   wire n1126;
   wire n1127;
   wire n1128;
   wire n1129;
   wire n1130;
   wire n1131;
   wire n1132;
   wire n1133;
   wire n1134;
   wire n1135;
   wire n1136;
   wire n1137;
   wire n1138;
   wire n1139;
   wire n1140;
   wire n1141;
   wire n1142;
   wire n1143;
   wire n1144;
   wire n1145;
   wire n1146;
   wire n1147;
   wire n1148;
   wire n1149;
   wire n1150;
   wire n1151;
   wire n1152;
   wire n1153;
   wire n1154;
   wire n1155;
   wire n1156;
   wire n1157;
   wire n1158;
   wire n1159;
   wire n1160;
   wire n1161;
   wire n1162;
   wire n1163;
   wire n1164;
   wire n1165;
   wire n1166;
   wire n1167;
   wire n1168;
   wire n1169;
   wire n1170;
   wire n1171;
   wire n1172;
   wire n1173;
   wire n1174;
   wire n1175;
   wire n1176;
   wire n1177;
   wire n1178;
   wire n1179;
   wire n1180;
   wire n1181;
   wire n1182;
   wire n1183;
   wire n1184;
   wire n1185;
   wire n1186;
   wire n1187;
   wire n1188;
   wire n1189;
   wire n1190;
   wire n1191;
   wire n1192;
   wire n1193;
   wire n1194;
   wire n1195;
   wire n1196;
   wire n1197;
   wire n1198;
   wire n1200;
   wire n1201;
   wire n1202;
   wire n1203;
   wire n1204;
   wire n1205;
   wire n1206;
   wire n1207;
   wire n1208;
   wire n1209;
   wire n1210;
   wire n1211;
   wire n1212;
   wire n1213;
   wire n1214;
   wire n1215;
   wire n1216;
   wire n1217;
   wire n1218;
   wire n1219;
   wire n1220;
   wire n1221;
   wire n1222;
   wire n1223;
   wire n1224;
   wire n1225;
   wire n1226;
   wire n1227;
   wire n1228;
   wire n1229;
   wire n1230;
   wire n1231;
   wire n1232;
   wire n1233;
   wire n1234;
   wire n1235;
   wire n1236;
   wire n1237;
   wire n1238;
   wire n1239;
   wire n1240;
   wire n1241;
   wire n1242;
   wire n1243;
   wire n1244;
   wire n1245;
   wire n1246;
   wire n1247;
   wire n1248;
   wire n1249;
   wire n1250;
   wire n1251;
   wire n1252;
   wire n1253;
   wire n1254;
   wire n1255;
   wire n1256;
   wire n1257;
   wire n1258;
   wire n1259;
   wire n1260;
   wire n1261;
   wire n1262;
   wire n1263;
   wire n1264;
   wire n1265;
   wire n1266;
   wire n1267;
   wire n1268;
   wire n1269;
   wire n1270;
   wire n1271;
   wire n1272;
   wire n1273;
   wire n1274;
   wire n1275;
   wire n1276;
   wire n1277;
   wire n1278;
   wire n1279;
   wire n1280;
   wire n1281;
   wire n1282;
   wire n1283;
   wire n1284;
   wire n1285;
   wire n1286;
   wire n1287;
   wire n1288;
   wire n1289;
   wire n1290;
   wire n1291;
   wire n1292;
   wire n1293;
   wire n1294;
   wire n1295;
   wire n1296;
   wire n1297;
   wire n1298;
   wire n1299;
   wire n1300;
   wire n1301;
   wire n1302;
   wire n1303;
   wire n1304;
   wire n1305;
   wire n1306;
   wire n1307;
   wire n1308;
   wire n1309;
   wire n1310;
   wire n1311;
   wire n1312;
   wire n1313;
   wire n1314;
   wire n1315;
   wire n1316;
   wire n1317;
   wire n1318;
   wire n1319;
   wire n1320;
   wire n1321;
   wire n1322;
   wire n1323;
   wire n1324;
   wire n1325;
   wire n1326;
   wire n1327;
   wire n1328;
   wire n1329;
   wire n1330;
   wire n1331;
   wire n1332;
   wire n1333;
   wire n1334;
   wire n1335;
   wire n1336;
   wire n1337;
   wire n1338;
   wire n1339;
   wire n1340;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n7;
   wire n8;
   wire n9;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n30;
   wire n35;
   wire n38;
   wire n39;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n83;
   wire n93;
   wire n96;
   wire n97;
   wire n99;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n110;
   wire n111;
   wire n113;
   wire n114;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n229;
   wire n705;
   wire n944;
   wire n1199;
   wire n1341;
   wire n1342;
   wire n1343;
   wire n1344;
   wire n1345;
   wire n1346;
   wire n1347;
   wire n1348;
   wire n1349;
   wire n1350;
   wire n1351;
   wire n1352;
   wire n1353;
   wire n1354;
   wire n1355;
   wire n1356;
   wire n1357;
   wire n1358;
   wire n1359;
   wire n1360;
   wire n1361;
   wire n1362;
   wire n1363;
   wire n1364;
   wire n1365;
   wire n1366;
   wire n1367;
   wire n1368;
   wire n1369;
   wire n1370;
   wire n1371;
   wire n1372;
   wire n1373;
   wire n1374;
   wire n1375;
   wire n1376;
   wire n1377;
   wire n1378;
   wire n1379;
   wire n1380;
   wire n1381;
   wire n1382;
   wire n1383;
   wire n1384;
   wire n1385;
   wire n1386;
   wire n1387;
   wire n1388;
   wire n1389;
   wire n1390;
   wire n1391;
   wire n1392;
   wire n1393;
   wire n1394;
   wire n1395;
   wire n1396;
   wire n1397;
   wire n1398;
   wire n1399;
   wire n1400;
   wire n1401;
   wire n1402;
   wire n1403;
   wire n1404;
   wire n1405;
   wire n1406;
   wire n1407;
   wire n1408;
   wire n1409;
   wire n1410;
   wire n1411;
   wire n1412;
   wire n1413;
   wire n1414;
   wire n1415;
   wire n1416;
   wire n1417;
   wire n1418;
   wire n1419;
   wire n1420;
   wire n1421;
   wire n1422;
   wire n1423;
   wire n1424;
   wire n1425;
   wire n1426;
   wire n1427;
   wire n1428;
   wire n1429;
   wire n1430;
   wire n1431;
   wire n1432;
   wire n1433;
   wire n1434;
   wire n1435;
   wire n1436;
   wire n1437;
   wire n1438;
   wire n1439;
   wire n1440;
   wire n1441;
   wire n1442;
   wire n1443;
   wire n1444;
   wire n1445;
   wire n1446;
   wire n1447;
   wire n1448;
   wire n1449;
   wire n1450;
   wire n1451;
   wire n1452;
   wire n1453;
   wire n1454;
   wire n1455;
   wire [1:0] sword_ctr_reg;
   wire [1:0] enc_ctrl_reg;

   BUFXL FE_PHC5256_n892 (.Y(FE_PHN5256_n892), 
	.A(n892));
   CLKBUFX1 FE_PHC5253_n1256 (.Y(FE_PHN5253_n1256), 
	.A(FE_PHN5227_n1256));
   BUFXL FE_PHC5252_n1296 (.Y(FE_PHN5252_n1296), 
	.A(FE_PHN5212_n1296));
   CLKBUFX1 FE_PHC5251_n866 (.Y(FE_PHN5251_n866), 
	.A(n866));
   BUFXL FE_PHC5250_n1264 (.Y(FE_PHN5250_n1264), 
	.A(FE_PHN5210_n1264));
   CLKBUFX1 FE_PHC5249_n1331 (.Y(FE_PHN5249_n1331), 
	.A(FE_PHN5211_n1331));
   BUFXL FE_PHC5248_n1236 (.Y(FE_PHN5248_n1236), 
	.A(FE_PHN5209_n1236));
   BUFXL FE_PHC5247_n1268 (.Y(FE_PHN5247_n1268), 
	.A(FE_PHN5199_n1268));
   BUFXL FE_PHC5246_n1276 (.Y(FE_PHN5246_n1276), 
	.A(FE_PHN5197_n1276));
   CLKBUFX1 FE_PHC5245_n1240 (.Y(FE_PHN5245_n1240), 
	.A(FE_PHN5208_n1240));
   CLKBUFX1 FE_PHC5244_n1138 (.Y(FE_PHN5244_n1138), 
	.A(FE_PHN5213_n1138));
   BUFXL FE_PHC5235_n658 (.Y(FE_PHN5235_n658), 
	.A(n658));
   CLKBUFX1 FE_PHC5233_n929 (.Y(FE_PHN5233_n929), 
	.A(n929));
   BUFXL FE_PHC5229_n1274 (.Y(FE_PHN5229_n1274), 
	.A(FE_PHN5117_n1274));
   CLKBUFX1 FE_PHC5228_n782 (.Y(FE_PHN5228_n782), 
	.A(n782));
   CLKBUFX1 FE_PHC5227_n1256 (.Y(FE_PHN5227_n1256), 
	.A(FE_PHN194_n1256));
   CLKBUFX1 FE_PHC5226_n1241 (.Y(FE_PHN5226_n1241), 
	.A(FE_PHN5108_n1241));
   DLY2X1 FE_PHC5225_n1238 (.Y(FE_PHN5225_n1238), 
	.A(n1238));
   BUFXL FE_PHC5224_n541 (.Y(FE_PHN5224_n541), 
	.A(n541));
   BUFXL FE_PHC5223_n1292 (.Y(FE_PHN5223_n1292), 
	.A(n1292));
   BUFXL FE_PHC5222_n1283 (.Y(FE_PHN5222_n1283), 
	.A(FE_PHN5151_n1283));
   BUFXL FE_PHC5221_n323 (.Y(FE_PHN5221_n323), 
	.A(n323));
   CLKBUFX1 FE_PHC5220_n1227 (.Y(FE_PHN5220_n1227), 
	.A(FE_PHN2805_n1227));
   CLKBUFX1 FE_PHC5219_n1252 (.Y(FE_PHN5219_n1252), 
	.A(FE_PHN241_n1252));
   CLKBUFX1 FE_PHC5218_n1279 (.Y(FE_PHN5218_n1279), 
	.A(FE_PHN196_n1279));
   CLKBUFX1 FE_PHC5217_n1266 (.Y(FE_PHN5217_n1266), 
	.A(FE_PHN5086_n1266));
   DLY2X1 FE_PHC5216_n1244 (.Y(FE_PHN5216_n1244), 
	.A(FE_PHN162_n1244));
   CLKBUFX1 FE_PHC5215_n1329 (.Y(FE_PHN5215_n1329), 
	.A(FE_PHN189_n1329));
   CLKBUFX1 FE_PHC5214_n774 (.Y(FE_PHN5214_n774), 
	.A(n774));
   BUFXL FE_PHC5213_n1138 (.Y(FE_PHN5213_n1138), 
	.A(n1138));
   CLKBUFX3 FE_PHC5212_n1296 (.Y(FE_PHN5212_n1296), 
	.A(n1296));
   CLKBUFX3 FE_PHC5211_n1331 (.Y(FE_PHN5211_n1331), 
	.A(FE_PHN188_n1331));
   CLKBUFX4 FE_PHC5210_n1264 (.Y(FE_PHN5210_n1264), 
	.A(FE_PHN158_n1264));
   CLKBUFX1 FE_PHC5209_n1236 (.Y(FE_PHN5209_n1236), 
	.A(FE_PHN182_n1236));
   BUFXL FE_PHC5208_n1240 (.Y(FE_PHN5208_n1240), 
	.A(FE_PHN5149_n1240));
   BUFXL FE_PHC5207_n866 (.Y(FE_PHN5207_n866), 
	.A(FE_PHN5251_n866));
   DLY2X1 FE_PHC5206_n316 (.Y(FE_PHN5206_n316), 
	.A(n316));
   BUFXL FE_PHC5205_n1273 (.Y(FE_PHN5205_n1273), 
	.A(n1273));
   DLY2X1 FE_PHC5204_n1229 (.Y(FE_PHN5204_n1229), 
	.A(n1229));
   DLY2X1 FE_PHC5203_n1209 (.Y(FE_PHN5203_n1209), 
	.A(n1209));
   DLY2X1 FE_PHC5202_n1272 (.Y(FE_PHN5202_n1272), 
	.A(FE_PHN118_n1272));
   DLY3X1 FE_PHC5201_n1225 (.Y(FE_PHN5201_n1225), 
	.A(FE_PHN183_n1225));
   BUFXL FE_PHC5200_n1249 (.Y(FE_PHN5200_n1249), 
	.A(n1249));
   CLKBUFX3 FE_PHC5199_n1268 (.Y(FE_PHN5199_n1268), 
	.A(n1268));
   DLY2X1 FE_PHC5198_n1208 (.Y(FE_PHN5198_n1208), 
	.A(n1208));
   CLKBUFX4 FE_PHC5197_n1276 (.Y(FE_PHN5197_n1276), 
	.A(FE_PHN5114_n1276));
   DLY2X1 FE_PHC5196_n1270 (.Y(FE_PHN5196_n1270), 
	.A(FE_PHN138_n1270));
   DLY2X1 FE_PHC5195_n1289 (.Y(FE_PHN5195_n1289), 
	.A(n1289));
   DLY2X1 FE_PHC5194_n1328 (.Y(FE_PHN5194_n1328), 
	.A(n1328));
   BUFXL FE_PHC5193_n1291 (.Y(FE_PHN5193_n1291), 
	.A(FE_PHN5092_n1291));
   DLY2X1 FE_PHC5192_n1265 (.Y(FE_PHN5192_n1265), 
	.A(FE_PHN5153_n1265));
   DLY2X1 FE_PHC5191_n1257 (.Y(FE_PHN5191_n1257), 
	.A(FE_PHN5141_n1257));
   DLY2X1 FE_PHC5190_n1280 (.Y(FE_PHN5190_n1280), 
	.A(n1280));
   DLY2X1 FE_PHC5189_n1248 (.Y(FE_PHN5189_n1248), 
	.A(n1248));
   DLY2X1 FE_PHC5188_n1218 (.Y(FE_PHN5188_n1218), 
	.A(n1218));
   DLY2X1 FE_PHC5187_n1233 (.Y(FE_PHN5187_n1233), 
	.A(FE_PHN5085_n1233));
   DLY1X1 FE_PHC5186_n1247 (.Y(FE_PHN5186_n1247), 
	.A(n1247));
   DLY2X1 FE_PHC5185_n1235 (.Y(FE_PHN5185_n1235), 
	.A(FE_PHN5080_n1235));
   DLY4X1 FE_PHC5184_n1219 (.Y(FE_PHN5184_n1219), 
	.A(FE_PHN5147_n1219));
   DLY2X1 FE_PHC5183_n1282 (.Y(FE_PHN5183_n1282), 
	.A(FE_PHN5098_n1282));
   DLY2X1 FE_PHC5182_n1242 (.Y(FE_PHN5182_n1242), 
	.A(FE_PHN5113_n1242));
   DLY2X1 FE_PHC5181_n1326 (.Y(FE_PHN5181_n1326), 
	.A(n1326));
   DLY3X1 FE_PHC5180_n1297 (.Y(FE_PHN5180_n1297), 
	.A(FE_PHN5104_n1297));
   DLY2X1 FE_PHC5179_n1269 (.Y(FE_PHN5179_n1269), 
	.A(FE_PHN5105_n1269));
   DLY2X1 FE_PHC5178_n1239 (.Y(FE_PHN5178_n1239), 
	.A(FE_PHN5139_n1239));
   DLY2X1 FE_PHC5177_n1324 (.Y(FE_PHN5177_n1324), 
	.A(FE_PHN5089_n1324));
   DLY3X1 FE_PHC5176_n1234 (.Y(FE_PHN5176_n1234), 
	.A(n1234));
   DLY2X1 FE_PHC5175_n1250 (.Y(FE_PHN5175_n1250), 
	.A(FE_PHN5138_n1250));
   DLY4X1 FE_PHC5174_n1232 (.Y(FE_PHN5174_n1232), 
	.A(n1232));
   BUFXL FE_PHC5172_n1100 (.Y(FE_PHN5172_n1100), 
	.A(n1100));
   BUFXL FE_PHC5169_n1297 (.Y(FE_PHN5169_n1297), 
	.A(FE_PHN5180_n1297));
   BUFXL FE_PHC5168_n1072 (.Y(FE_PHN5168_n1072), 
	.A(FE_PHN5137_n1072));
   BUFXL FE_PHC5167_n1028 (.Y(FE_PHN5167_n1028), 
	.A(FE_PHN5112_n1028));
   CLKBUFX1 FE_PHC5166_n1219 (.Y(FE_PHN5166_n1219), 
	.A(FE_PHN5184_n1219));
   BUFXL FE_PHC5165_n563 (.Y(FE_PHN5165_n563), 
	.A(FE_PHN5103_n563));
   CLKBUFX1 FE_PHC5164_n1131 (.Y(FE_PHN5164_n1131), 
	.A(n1131));
   CLKBUFX1 FE_PHC5163_n1291 (.Y(FE_PHN5163_n1291), 
	.A(FE_PHN5193_n1291));
   CLKBUFX1 FE_PHC5162_n1274 (.Y(FE_PHN5162_n1274), 
	.A(FE_PHN5229_n1274));
   BUFXL FE_PHC5161_n426 (.Y(FE_PHN5161_n426), 
	.A(FE_PHN5128_n426));
   CLKBUFX1 FE_PHC5160_n1307 (.Y(FE_PHN5160_n1307), 
	.A(FE_PHN5129_n1307));
   BUFXL FE_PHC5153_n1265 (.Y(FE_PHN5153_n1265), 
	.A(FE_PHN159_n1265));
   BUFXL FE_PHC5152_n1090 (.Y(FE_PHN5152_n1090), 
	.A(n1090));
   BUFXL FE_PHC5151_n1283 (.Y(FE_PHN5151_n1283), 
	.A(n1283));
   BUFXL FE_PHC5150_n782 (.Y(FE_PHN5150_n782), 
	.A(FE_PHN5228_n782));
   CLKBUFX1 FE_PHC5149_n1240 (.Y(FE_PHN5149_n1240), 
	.A(n1240));
   CLKBUFX1 FE_PHC5148_n372 (.Y(FE_PHN5148_n372), 
	.A(n372));
   CLKBUFX3 FE_PHC5147_n1219 (.Y(FE_PHN5147_n1219), 
	.A(n1219));
   CLKBUFX1 FE_PHC5146_n548 (.Y(FE_PHN5146_n548), 
	.A(n548));
   BUFXL FE_PHC5145_n1302 (.Y(FE_PHN5145_n1302), 
	.A(FE_PHN143_n1302));
   CLKBUFX1 FE_PHC5144_n1078 (.Y(FE_PHN5144_n1078), 
	.A(n1078));
   BUFXL FE_PHC5143_n1305 (.Y(FE_PHN5143_n1305), 
	.A(FE_PHN125_n1305));
   BUFXL FE_PHC5142_n309 (.Y(FE_PHN5142_n309), 
	.A(n309));
   BUFXL FE_PHC5141_n1257 (.Y(FE_PHN5141_n1257), 
	.A(n1257));
   BUFXL FE_PHC5140_n1206 (.Y(FE_PHN5140_n1206), 
	.A(n1206));
   BUFXL FE_PHC5139_n1239 (.Y(FE_PHN5139_n1239), 
	.A(n1239));
   CLKBUFX1 FE_PHC5138_n1250 (.Y(FE_PHN5138_n1250), 
	.A(n1250));
   CLKBUFX1 FE_PHC5137_n1072 (.Y(FE_PHN5137_n1072), 
	.A(n1072));
   DLY2X1 FE_PHC5136_n1251 (.Y(FE_PHN5136_n1251), 
	.A(FE_PHN174_n1251));
   BUFXL FE_PHC5135_n1237 (.Y(FE_PHN5135_n1237), 
	.A(n1237));
   BUFXL FE_PHC5134_n541 (.Y(FE_PHN5134_n541), 
	.A(FE_PHN5224_n541));
   DLY1X1 FE_PHC5133_n1043 (.Y(FE_PHN5133_n1043), 
	.A(n1043));
   DLY2X1 FE_PHC5132_n378 (.Y(FE_PHN5132_n378), 
	.A(n378));
   DLY2X1 FE_PHC5131_n1300 (.Y(FE_PHN5131_n1300), 
	.A(n1300));
   CLKBUFX1 FE_PHC5130_n1210 (.Y(FE_PHN5130_n1210), 
	.A(n1210));
   CLKBUFX3 FE_PHC5129_n1307 (.Y(FE_PHN5129_n1307), 
	.A(n1307));
   CLKBUFX3 FE_PHC5128_n426 (.Y(FE_PHN5128_n426), 
	.A(n426));
   CLKBUFX1 FE_PHC5127_n1035 (.Y(FE_PHN5127_n1035), 
	.A(n1035));
   CLKBUFX1 FE_PHC5126_n1021 (.Y(FE_PHN5126_n1021), 
	.A(n1021));
   DLY2X1 FE_PHC5125_n366 (.Y(FE_PHN5125_n366), 
	.A(n366));
   DLY2X1 FE_PHC5124_n1212 (.Y(FE_PHN5124_n1212), 
	.A(n1212));
   DLY2X1 FE_PHC5123_n1323 (.Y(FE_PHN5123_n1323), 
	.A(n1323));
   DLY2X1 FE_PHC5122_n1213 (.Y(FE_PHN5122_n1213), 
	.A(n1213));
   DLY2X1 FE_PHC5121_n1314 (.Y(FE_PHN5121_n1314), 
	.A(FE_PHN210_n1314));
   BUFXL FE_PHC5120_n1230 (.Y(FE_PHN5120_n1230), 
	.A(n1230));
   CLKBUFX1 FE_PHC5119_n651 (.Y(FE_PHN5119_n651), 
	.A(n651));
   CLKBUFX1 FE_PHC5118_n1308 (.Y(FE_PHN5118_n1308), 
	.A(n1308));
   CLKBUFX1 FE_PHC5117_n1274 (.Y(FE_PHN5117_n1274), 
	.A(n1274));
   DLY2X1 FE_PHC5116_n1322 (.Y(FE_PHN5116_n1322), 
	.A(n1322));
   CLKBUFX1 FE_PHC5115_n1303 (.Y(FE_PHN5115_n1303), 
	.A(n1303));
   CLKBUFX1 FE_PHC5114_n1276 (.Y(FE_PHN5114_n1276), 
	.A(n1276));
   CLKBUFX1 FE_PHC5113_n1242 (.Y(FE_PHN5113_n1242), 
	.A(n1242));
   CLKBUFX1 FE_PHC5112_n1028 (.Y(FE_PHN5112_n1028), 
	.A(n1028));
   DLY2X1 FE_PHC5111_n1275 (.Y(FE_PHN5111_n1275), 
	.A(FE_PHN128_n1275));
   DLY2X1 FE_PHC5110_n441 (.Y(FE_PHN5110_n441), 
	.A(n441));
   DLY2X1 FE_PHC5109_n696 (.Y(FE_PHN5109_n696), 
	.A(n696));
   DLY2X1 FE_PHC5108_n1241 (.Y(FE_PHN5108_n1241), 
	.A(FE_PHN133_n1241));
   DLY2X1 FE_PHC5107_n1220 (.Y(FE_PHN5107_n1220), 
	.A(FE_PHN177_n1220));
   DLY2X1 FE_PHC5106_n1315 (.Y(FE_PHN5106_n1315), 
	.A(FE_PHN176_n1315));
   CLKBUFX1 FE_PHC5105_n1269 (.Y(FE_PHN5105_n1269), 
	.A(n1269));
   CLKBUFX1 FE_PHC5104_n1297 (.Y(FE_PHN5104_n1297), 
	.A(n1297));
   CLKBUFX1 FE_PHC5103_n563 (.Y(FE_PHN5103_n563), 
	.A(n563));
   BUFXL FE_PHC5102_n1131 (.Y(FE_PHN5102_n1131), 
	.A(FE_PHN5164_n1131));
   DLY2X1 FE_PHC5101_n1066 (.Y(FE_PHN5101_n1066), 
	.A(n1066));
   DLY2X1 FE_PHC5100_n1244 (.Y(FE_PHN5100_n1244), 
	.A(n1244));
   DLY2X1 FE_PHC5099_n1243 (.Y(FE_PHN5099_n1243), 
	.A(n1243));
   CLKBUFX1 FE_PHC5098_n1282 (.Y(FE_PHN5098_n1282), 
	.A(FE_PHN205_n1282));
   DLY2X1 FE_PHC5097_n1333 (.Y(FE_PHN5097_n1333), 
	.A(FE_PHN206_n1333));
   DLY2X1 FE_PHC5096_n1221 (.Y(FE_PHN5096_n1221), 
	.A(FE_PHN252_n1221));
   DLY2X1 FE_PHC5095_n1211 (.Y(FE_PHN5095_n1211), 
	.A(FE_PHN134_n1211));
   DLY2X1 FE_PHC5094_n1267 (.Y(FE_PHN5094_n1267), 
	.A(n1267));
   DLY2X1 FE_PHC5093_n1236 (.Y(FE_PHN5093_n1236), 
	.A(n1236));
   CLKBUFX3 FE_PHC5092_n1291 (.Y(FE_PHN5092_n1291), 
	.A(n1291));
   DLY2X1 FE_PHC5091_n1098 (.Y(FE_PHN5091_n1098), 
	.A(n1098));
   DLY2X1 FE_PHC5090_n1306 (.Y(FE_PHN5090_n1306), 
	.A(n1306));
   DLY2X1 FE_PHC5089_n1324 (.Y(FE_PHN5089_n1324), 
	.A(FE_PHN245_n1324));
   DLY2X1 FE_PHC5088_n1281 (.Y(FE_PHN5088_n1281), 
	.A(n1281));
   DLY2X1 FE_PHC5087_n1304 (.Y(FE_PHN5087_n1304), 
	.A(n1304));
   DLY2X1 FE_PHC5086_n1266 (.Y(FE_PHN5086_n1266), 
	.A(FE_PHN181_n1266));
   DLY2X1 FE_PHC5085_n1233 (.Y(FE_PHN5085_n1233), 
	.A(FE_PHN164_n1233));
   DLY2X1 FE_PHC5084_n1226 (.Y(FE_PHN5084_n1226), 
	.A(n1226));
   DLY2X1 FE_PHC5083_n1228 (.Y(FE_PHN5083_n1228), 
	.A(n1228));
   DLY4X1 FE_PHC5082_n1245 (.Y(FE_PHN5082_n1245), 
	.A(n1245));
   DLY1X1 FE_PHC5081_n1290 (.Y(FE_PHN5081_n1290), 
	.A(FE_PHN230_n1290));
   DLY2X1 FE_PHC5080_n1235 (.Y(FE_PHN5080_n1235), 
	.A(FE_PHN204_n1235));
   DLY2X1 FE_PHC5079_n1299 (.Y(FE_PHN5079_n1299), 
	.A(FE_PHN167_n1299));
   DLY2X1 FE_PHC5078_n1258 (.Y(FE_PHN5078_n1258), 
	.A(n1258));
   BUFXL FE_PHC5075_n419 (.Y(FE_PHN5075_n419), 
	.A(n419));
   DLY2X1 FE_PHC5045_n1334 (.Y(FE_PHN5045_n1334), 
	.A(n1334));
   DLY4X1 FE_PHC3408_enc_ctrl_reg_0_ (.Y(FE_PHN3408_enc_ctrl_reg_0_), 
	.A(FE_PHN410_enc_ctrl_reg_0_));
   DLY4X1 FE_PHC3108_Dout_104_ (.Y(new_block[104]), 
	.A(FE_PHN3108_Dout_104_));
   DLY3X1 FE_PHC3107_Dout_33_ (.Y(new_block[33]), 
	.A(FE_PHN3107_Dout_33_));
   DLY4X1 FE_PHC3106_Dout_97_ (.Y(new_block[97]), 
	.A(FE_PHN3106_Dout_97_));
   DLY3X1 FE_PHC3105_Dout_47_ (.Y(new_block[47]), 
	.A(FE_PHN3105_Dout_47_));
   DLY4X1 FE_PHC3104_Dout_8_ (.Y(new_block[8]), 
	.A(FE_PHN3104_Dout_8_));
   DLY3X1 FE_PHC3095_Dout_119_ (.Y(new_block[119]), 
	.A(FE_PHN3095_Dout_119_));
   DLY2X1 FE_PHC3081_n1194 (.Y(FE_PHN3081_n1194), 
	.A(n1194));
   DLY2X1 FE_PHC2856_n1338 (.Y(FE_PHN2856_n1338), 
	.A(n1338));
   DLY2X1 FE_PHC2850_Dout_125_ (.Y(new_block[125]), 
	.A(FE_PHN2850_Dout_125_));
   DLY2X1 FE_PHC2843_n1335 (.Y(FE_PHN2843_n1335), 
	.A(n1335));
   DLY2X1 FE_PHC2821_enc_ctrl_reg_1_ (.Y(FE_PHN2821_enc_ctrl_reg_1_), 
	.A(FE_PHN111_enc_ctrl_reg_1_));
   DLY4X1 FE_PHC2816_n1013 (.Y(FE_PHN2816_n1013), 
	.A(n1013));
   DLY2X1 FE_PHC2813_enc_round_nr_2_ (.Y(FE_PHN2813_enc_round_nr_2_), 
	.A(round[2]));
   DLY2X1 FE_PHC2812_enc_round_nr_1_ (.Y(round[1]), 
	.A(FE_PHN2812_enc_round_nr_1_));
   DLY4X1 FE_PHC2809_n1340 (.Y(FE_PHN2809_n1340), 
	.A(n1340));
   CLKBUFX3 FE_PHC2807_n1330 (.Y(FE_PHN2807_n1330), 
	.A(FE_PHN213_n1330));
   DLY2X1 FE_PHC2806_n1301 (.Y(FE_PHN2806_n1301), 
	.A(n1301));
   DLY1X1 FE_PHC2805_n1227 (.Y(FE_PHN2805_n1227), 
	.A(n1227));
   DLY4X1 FE_PHC1310_n1334 (.Y(FE_PHN1310_n1334), 
	.A(FE_PHN5045_n1334));
   DLY4X1 FE_PHC821_Dout_1_ (.Y(new_block[1]), 
	.A(FE_PHN821_Dout_1_));
   DLY4X1 FE_PHC751_n1337 (.Y(FE_PHN751_n1337), 
	.A(n1337));
   DLY4X1 FE_PHC750_Dout_103_ (.Y(new_block[103]), 
	.A(FE_PHN750_Dout_103_));
   DLY4X1 FE_PHC703_n1336 (.Y(FE_PHN703_n1336), 
	.A(n1336));
   DLY4X1 FE_PHC702_Dout_38_ (.Y(new_block[38]), 
	.A(FE_PHN702_Dout_38_));
   DLY4X1 FE_PHC701_Dout_36_ (.Y(new_block[36]), 
	.A(FE_PHN701_Dout_36_));
   DLY4X1 FE_PHC604_Dout_34_ (.Y(new_block[34]), 
	.A(FE_PHN604_Dout_34_));
   DLY4X1 FE_PHC603_Dout_10_ (.Y(new_block[10]), 
	.A(FE_PHN603_Dout_10_));
   DLY4X1 FE_PHC602_n1197 (.Y(FE_PHN602_n1197), 
	.A(n1197));
   DLY4X1 FE_PHC601_Dout_46_ (.Y(new_block[46]), 
	.A(FE_PHN601_Dout_46_));
   DLY4X1 FE_PHC600_Dout_37_ (.Y(new_block[37]), 
	.A(FE_PHN600_Dout_37_));
   DLY4X1 FE_PHC599_Dout_102_ (.Y(new_block[102]), 
	.A(FE_PHN599_Dout_102_));
   DLY4X1 FE_PHC598_Dout_116_ (.Y(new_block[116]), 
	.A(FE_PHN598_Dout_116_));
   DLY4X1 FE_PHC597_Dout_44_ (.Y(new_block[44]), 
	.A(FE_PHN597_Dout_44_));
   DLY4X1 FE_PHC596_Dout_101_ (.Y(new_block[101]), 
	.A(FE_PHN596_Dout_101_));
   DLY4X1 FE_PHC595_Dout_110_ (.Y(new_block[110]), 
	.A(FE_PHN595_Dout_110_));
   DLY4X1 FE_PHC535_enc_ctrl_we (.Y(FE_PHN535_enc_ctrl_we), 
	.A(enc_ctrl_we));
   DLY4X1 FE_PHC533_Dout_122_ (.Y(new_block[122]), 
	.A(FE_PHN533_Dout_122_));
   DLY4X1 FE_PHC528_Dout_111_ (.Y(new_block[111]), 
	.A(FE_PHN528_Dout_111_));
   DLY4X1 FE_PHC444_Dout_73_ (.Y(new_block[73]), 
	.A(FE_PHN444_Dout_73_));
   DLY4X1 FE_PHC443_Dout_72_ (.Y(new_block[72]), 
	.A(FE_PHN443_Dout_72_));
   DLY4X1 FE_PHC442_Dout_114_ (.Y(new_block[114]), 
	.A(FE_PHN442_Dout_114_));
   DLY4X1 FE_PHC441_Dout_9_ (.Y(new_block[9]), 
	.A(FE_PHN441_Dout_9_));
   DLY4X1 FE_PHC440_Dout_54_ (.Y(new_block[54]), 
	.A(FE_PHN440_Dout_54_));
   DLY4X1 FE_PHC438_Dout_0_ (.Y(new_block[0]), 
	.A(FE_PHN438_Dout_0_));
   DLY4X1 FE_PHC437_Dout_108_ (.Y(new_block[108]), 
	.A(FE_PHN437_Dout_108_));
   DLY4X1 FE_PHC436_Dout_117_ (.Y(new_block[117]), 
	.A(FE_PHN436_Dout_117_));
   DLY4X1 FE_PHC435_Dout_109_ (.Y(new_block[109]), 
	.A(FE_PHN435_Dout_109_));
   DLY4X1 FE_PHC433_Dout_100_ (.Y(new_block[100]), 
	.A(FE_PHN433_Dout_100_));
   DLY4X1 FE_PHC415_Dout_93_ (.Y(new_block[93]), 
	.A(FE_PHN415_Dout_93_));
   DLY4X1 FE_PHC414_Dout_63_ (.Y(new_block[63]), 
	.A(FE_PHN414_Dout_63_));
   DLY4X1 FE_PHC413_Dout_120_ (.Y(new_block[120]), 
	.A(FE_PHN413_Dout_120_));
   DLY4X1 FE_PHC412_Dout_126_ (.Y(new_block[126]), 
	.A(FE_PHN412_Dout_126_));
   DLY4X1 FE_PHC410_enc_ctrl_reg_0_ (.Y(FE_PHN410_enc_ctrl_reg_0_), 
	.A(enc_ctrl_reg[0]));
   DLY4X1 FE_PHC378_Dout_39_ (.Y(new_block[39]), 
	.A(FE_PHN378_Dout_39_));
   DLY4X1 FE_PHC377_Dout_6_ (.Y(new_block[6]), 
	.A(FE_PHN377_Dout_6_));
   DLY4X1 FE_PHC374_Dout_53_ (.Y(new_block[53]), 
	.A(FE_PHN374_Dout_53_));
   DLY4X1 FE_PHC373_Dout_68_ (.Y(new_block[68]), 
	.A(FE_PHN373_Dout_68_));
   DLY4X1 FE_PHC371_Dout_35_ (.Y(new_block[35]), 
	.A(FE_PHN371_Dout_35_));
   DLY4X1 FE_PHC369_Dout_105_ (.Y(new_block[105]), 
	.A(FE_PHN369_Dout_105_));
   DLY4X1 FE_PHC368_Dout_74_ (.Y(new_block[74]), 
	.A(FE_PHN368_Dout_74_));
   DLY4X1 FE_PHC367_Dout_76_ (.Y(new_block[76]), 
	.A(FE_PHN367_Dout_76_));
   DLY4X1 FE_PHC366_Dout_20_ (.Y(new_block[20]), 
	.A(FE_PHN366_Dout_20_));
   DLY4X1 FE_PHC365_Dout_22_ (.Y(new_block[22]), 
	.A(FE_PHN365_Dout_22_));
   DLY4X1 FE_PHC364_Dout_21_ (.Y(new_block[21]), 
	.A(FE_PHN364_Dout_21_));
   DLY4X1 FE_PHC363_Dout_3_ (.Y(new_block[3]), 
	.A(FE_PHN363_Dout_3_));
   DLY4X1 FE_PHC362_Dout_45_ (.Y(new_block[45]), 
	.A(FE_PHN362_Dout_45_));
   DLY4X1 FE_PHC361_Dout_127_ (.Y(new_block[127]), 
	.A(FE_PHN361_Dout_127_));
   DLY4X1 FE_PHC356_Dout_26_ (.Y(new_block[26]), 
	.A(FE_PHN356_Dout_26_));
   DLY4X1 FE_PHC355_Dout_58_ (.Y(new_block[58]), 
	.A(FE_PHN355_Dout_58_));
   DLY4X1 FE_PHC354_n1335 (.Y(FE_PHN354_n1335), 
	.A(FE_PHN2843_n1335));
   DLY4X1 FE_PHC353_Dout_60_ (.Y(new_block[60]), 
	.A(FE_PHN353_Dout_60_));
   DLY4X1 FE_PHC352_Dout_123_ (.Y(new_block[123]), 
	.A(FE_PHN352_Dout_123_));
   DLY4X1 FE_PHC351_Dout_121_ (.Y(new_block[121]), 
	.A(FE_PHN351_Dout_121_));
   DLY4X1 FE_PHC350_Dout_124_ (.Y(new_block[124]), 
	.A(FE_PHN350_Dout_124_));
   DLY4X1 FE_PHC341_Dout_79_ (.Y(new_block[79]), 
	.A(FE_PHN341_Dout_79_));
   DLY4X1 FE_PHC340_Dout_65_ (.Y(new_block[65]), 
	.A(FE_PHN340_Dout_65_));
   DLY4X1 FE_PHC339_Dout_107_ (.Y(new_block[107]), 
	.A(FE_PHN339_Dout_107_));
   DLY4X1 FE_PHC338_Dout_11_ (.Y(new_block[11]), 
	.A(FE_PHN338_Dout_11_));
   DLY4X1 FE_PHC337_Dout_115_ (.Y(new_block[115]), 
	.A(FE_PHN337_Dout_115_));
   DLY4X1 FE_PHC336_Dout_15_ (.Y(new_block[15]), 
	.A(FE_PHN336_Dout_15_));
   DLY4X1 FE_PHC335_Dout_112_ (.Y(new_block[112]), 
	.A(FE_PHN335_Dout_112_));
   DLY4X1 FE_PHC334_Dout_49_ (.Y(new_block[49]), 
	.A(FE_PHN334_Dout_49_));
   DLY4X1 FE_PHC333_Dout_48_ (.Y(new_block[48]), 
	.A(FE_PHN333_Dout_48_));
   DLY4X1 FE_PHC332_Dout_52_ (.Y(new_block[52]), 
	.A(FE_PHN332_Dout_52_));
   DLY4X1 FE_PHC331_Dout_17_ (.Y(new_block[17]), 
	.A(FE_PHN331_Dout_17_));
   DLY4X1 FE_PHC330_Dout_118_ (.Y(new_block[118]), 
	.A(FE_PHN330_Dout_118_));
   DLY4X1 FE_PHC329_Dout_4_ (.Y(new_block[4]), 
	.A(FE_PHN329_Dout_4_));
   DLY4X1 FE_PHC328_Dout_113_ (.Y(new_block[113]), 
	.A(FE_PHN328_Dout_113_));
   DLY4X1 FE_PHC321_Dout_90_ (.Y(new_block[90]), 
	.A(FE_PHN321_Dout_90_));
   DLY4X1 FE_PHC320_Dout_88_ (.Y(new_block[88]), 
	.A(FE_PHN320_Dout_88_));
   DLY4X1 FE_PHC318_Dout_62_ (.Y(new_block[62]), 
	.A(FE_PHN318_Dout_62_));
   DLY4X1 FE_PHC317_Dout_19_ (.Y(new_block[19]), 
	.A(FE_PHN317_Dout_19_));
   DLY4X1 FE_PHC316_Dout_85_ (.Y(new_block[85]), 
	.A(FE_PHN316_Dout_85_));
   DLY4X1 FE_PHC315_Dout_42_ (.Y(new_block[42]), 
	.A(FE_PHN315_Dout_42_));
   DLY4X1 FE_PHC314_Dout_18_ (.Y(new_block[18]), 
	.A(FE_PHN314_Dout_18_));
   DLY4X1 FE_PHC313_Dout_32_ (.Y(new_block[32]), 
	.A(FE_PHN313_Dout_32_));
   DLY4X1 FE_PHC312_Dout_50_ (.Y(new_block[50]), 
	.A(FE_PHN312_Dout_50_));
   DLY4X1 FE_PHC311_Dout_99_ (.Y(new_block[99]), 
	.A(FE_PHN311_Dout_99_));
   DLY4X1 FE_PHC310_Dout_16_ (.Y(new_block[16]), 
	.A(FE_PHN310_Dout_16_));
   DLY4X1 FE_PHC309_Dout_70_ (.Y(new_block[70]), 
	.A(FE_PHN309_Dout_70_));
   DLY4X1 FE_PHC308_Dout_80_ (.Y(new_block[80]), 
	.A(FE_PHN308_Dout_80_));
   DLY4X1 FE_PHC307_Dout_13_ (.Y(new_block[13]), 
	.A(FE_PHN307_Dout_13_));
   DLY4X1 FE_PHC306_Dout_51_ (.Y(new_block[51]), 
	.A(FE_PHN306_Dout_51_));
   DLY4X1 FE_PHC305_Dout_41_ (.Y(new_block[41]), 
	.A(FE_PHN305_Dout_41_));
   DLY4X1 FE_PHC304_Dout_95_ (.Y(new_block[95]), 
	.A(FE_PHN304_Dout_95_));
   DLY4X1 FE_PHC303_Dout_92_ (.Y(new_block[92]), 
	.A(FE_PHN303_Dout_92_));
   DLY4X1 FE_PHC302_Dout_28_ (.Y(new_block[28]), 
	.A(FE_PHN302_Dout_28_));
   DLY4X1 FE_PHC300_Dout_55_ (.Y(new_block[55]), 
	.A(FE_PHN300_Dout_55_));
   DLY4X1 FE_PHC299_Dout_23_ (.Y(new_block[23]), 
	.A(FE_PHN299_Dout_23_));
   DLY4X1 FE_PHC298_Dout_7_ (.Y(new_block[7]), 
	.A(FE_PHN298_Dout_7_));
   DLY4X1 FE_PHC297_Dout_64_ (.Y(new_block[64]), 
	.A(FE_PHN297_Dout_64_));
   DLY4X1 FE_PHC296_Dout_84_ (.Y(new_block[84]), 
	.A(FE_PHN296_Dout_84_));
   DLY4X1 FE_PHC295_Dout_14_ (.Y(new_block[14]), 
	.A(FE_PHN295_Dout_14_));
   DLY4X1 FE_PHC294_Dout_77_ (.Y(new_block[77]), 
	.A(FE_PHN294_Dout_77_));
   DLY4X1 FE_PHC293_Dout_75_ (.Y(new_block[75]), 
	.A(FE_PHN293_Dout_75_));
   DLY4X1 FE_PHC292_Dout_78_ (.Y(new_block[78]), 
	.A(FE_PHN292_Dout_78_));
   DLY4X1 FE_PHC289_Dout_91_ (.Y(new_block[91]), 
	.A(FE_PHN289_Dout_91_));
   DLY4X1 FE_PHC288_Dout_94_ (.Y(new_block[94]), 
	.A(FE_PHN288_Dout_94_));
   DLY4X1 FE_PHC287_Dout_59_ (.Y(new_block[59]), 
	.A(FE_PHN287_Dout_59_));
   DLY4X1 FE_PHC286_Dout_24_ (.Y(new_block[24]), 
	.A(FE_PHN286_Dout_24_));
   DLY4X1 FE_PHC285_Dout_25_ (.Y(new_block[25]), 
	.A(FE_PHN285_Dout_25_));
   DLY4X1 FE_PHC284_Dout_57_ (.Y(new_block[57]), 
	.A(FE_PHN284_Dout_57_));
   DLY4X1 FE_PHC282_Dout_30_ (.Y(new_block[30]), 
	.A(FE_PHN282_Dout_30_));
   DLY4X1 FE_PHC281_Dout_31_ (.Y(new_block[31]), 
	.A(FE_PHN281_Dout_31_));
   DLY4X1 FE_PHC280_Dout_40_ (.Y(new_block[40]), 
	.A(FE_PHN280_Dout_40_));
   DLY4X1 FE_PHC279_Dout_86_ (.Y(new_block[86]), 
	.A(FE_PHN279_Dout_86_));
   DLY4X1 FE_PHC278_Dout_87_ (.Y(new_block[87]), 
	.A(FE_PHN278_Dout_87_));
   DLY4X1 FE_PHC277_Dout_81_ (.Y(new_block[81]), 
	.A(FE_PHN277_Dout_81_));
   DLY4X1 FE_PHC276_Dout_67_ (.Y(new_block[67]), 
	.A(FE_PHN276_Dout_67_));
   DLY4X1 FE_PHC275_Dout_12_ (.Y(new_block[12]), 
	.A(FE_PHN275_Dout_12_));
   DLY4X1 FE_PHC274_Dout_82_ (.Y(new_block[82]), 
	.A(FE_PHN274_Dout_82_));
   DLY4X1 FE_PHC273_Dout_66_ (.Y(new_block[66]), 
	.A(FE_PHN273_Dout_66_));
   DLY4X1 FE_PHC272_Dout_89_ (.Y(new_block[89]), 
	.A(FE_PHN272_Dout_89_));
   DLY4X1 FE_PHC269_Dout_71_ (.Y(new_block[71]), 
	.A(FE_PHN269_Dout_71_));
   DLY4X1 FE_PHC268_Dout_96_ (.Y(new_block[96]), 
	.A(FE_PHN268_Dout_96_));
   DLY4X1 FE_PHC267_Dout_83_ (.Y(new_block[83]), 
	.A(FE_PHN267_Dout_83_));
   DLY4X1 FE_PHC266_Dout_98_ (.Y(new_block[98]), 
	.A(FE_PHN266_Dout_98_));
   DLY4X1 FE_PHC264_Dout_27_ (.Y(new_block[27]), 
	.A(FE_PHN264_Dout_27_));
   DLY4X1 FE_PHC263_Dout_56_ (.Y(new_block[56]), 
	.A(FE_PHN263_Dout_56_));
   DLY4X1 FE_PHC262_Dout_61_ (.Y(new_block[61]), 
	.A(FE_PHN262_Dout_61_));
   DLY4X1 FE_PHC261_Dout_69_ (.Y(new_block[69]), 
	.A(FE_PHN261_Dout_69_));
   DLY4X1 FE_PHC260_Dout_43_ (.Y(new_block[43]), 
	.A(FE_PHN260_Dout_43_));
   DLY4X1 FE_PHC259_Dout_5_ (.Y(new_block[5]), 
	.A(FE_PHN259_Dout_5_));
   DLY4X1 FE_PHC258_n1339 (.Y(FE_PHN258_n1339), 
	.A(n1339));
   DLY4X1 FE_PHC257_Dout_29_ (.Y(new_block[29]), 
	.A(FE_PHN257_Dout_29_));
   DLY4X1 FE_PHC256_n943 (.Y(FE_PHN256_n943), 
	.A(n943));
   DLY4X1 FE_PHC253_n704 (.Y(FE_PHN253_n704), 
	.A(n704));
   DLY4X1 FE_PHC252_n1221 (.Y(FE_PHN252_n1221), 
	.A(n1221));
   DLY4X1 FE_PHC251_n1229 (.Y(FE_PHN251_n1229), 
	.A(FE_PHN5204_n1229));
   DLY4X1 FE_PHC250_n1223 (.Y(FE_PHN250_n1223), 
	.A(n1223));
   DLY4X1 FE_PHC249_n1222 (.Y(FE_PHN249_n1222), 
	.A(n1222));
   DLY4X1 FE_PHC248_n1316 (.Y(FE_PHN248_n1316), 
	.A(n1316));
   DLY4X1 FE_PHC247_n1332 (.Y(FE_PHN247_n1332), 
	.A(n1332));
   DLY4X1 FE_PHC246_n1317 (.Y(FE_PHN246_n1317), 
	.A(n1317));
   DLY4X1 FE_PHC245_n1324 (.Y(FE_PHN245_n1324), 
	.A(n1324));
   DLY4X1 FE_PHC244_n1322 (.Y(FE_PHN244_n1322), 
	.A(FE_PHN5116_n1322));
   DLY4X1 FE_PHC243_n1224 (.Y(FE_PHN243_n1224), 
	.A(n1224));
   DLY4X1 FE_PHC242_n1318 (.Y(FE_PHN242_n1318), 
	.A(n1318));
   DLY4X1 FE_PHC241_n1252 (.Y(FE_PHN241_n1252), 
	.A(n1252));
   DLY4X1 FE_PHC240_n1287 (.Y(FE_PHN240_n1287), 
	.A(n1287));
   DLY4X1 FE_PHC239_n1284 (.Y(FE_PHN239_n1284), 
	.A(n1284));
   DLY4X1 FE_PHC238_n1319 (.Y(FE_PHN238_n1319), 
	.A(n1319));
   DLY4X1 FE_PHC237_n1254 (.Y(FE_PHN237_n1254), 
	.A(n1254));
   DLY4X1 FE_PHC236_n1292 (.Y(FE_PHN236_n1292), 
	.A(FE_PHN5223_n1292));
   DLY4X1 FE_PHC235_n1285 (.Y(FE_PHN235_n1285), 
	.A(n1285));
   DLY4X1 FE_PHC234_n1255 (.Y(FE_PHN234_n1255), 
	.A(n1255));
   DLY4X1 FE_PHC233_n1253 (.Y(FE_PHN233_n1253), 
	.A(n1253));
   DLY4X1 FE_PHC232_n1286 (.Y(FE_PHN232_n1286), 
	.A(n1286));
   DLY4X1 FE_PHC231_n1227 (.Y(FE_PHN231_n1227), 
	.A(FE_PHN5220_n1227));
   DLY4X1 FE_PHC230_n1290 (.Y(FE_PHN230_n1290), 
	.A(n1290));
   DLY4X1 FE_PHC229_n1216 (.Y(FE_PHN229_n1216), 
	.A(n1216));
   DLY4X1 FE_PHC228_n1300 (.Y(FE_PHN228_n1300), 
	.A(FE_PHN5131_n1300));
   DLY4X1 FE_PHC227_n1258 (.Y(FE_PHN227_n1258), 
	.A(FE_PHN5078_n1258));
   DLY4X1 FE_PHC226_n1214 (.Y(FE_PHN226_n1214), 
	.A(n1214));
   DLY4X1 FE_PHC225_n1277 (.Y(FE_PHN225_n1277), 
	.A(n1277));
   DLY4X1 FE_PHC224_n1327 (.Y(FE_PHN224_n1327), 
	.A(n1327));
   DLY4X1 FE_PHC223_n1228 (.Y(FE_PHN223_n1228), 
	.A(FE_PHN5083_n1228));
   DLY4X1 FE_PHC222_n1215 (.Y(FE_PHN222_n1215), 
	.A(n1215));
   DLY4X1 FE_PHC221_n1309 (.Y(FE_PHN221_n1309), 
	.A(n1309));
   DLY4X1 FE_PHC220_n1311 (.Y(FE_PHN220_n1311), 
	.A(n1311));
   DLY4X1 FE_PHC219_n1232 (.Y(FE_PHN219_n1232), 
	.A(FE_PHN5174_n1232));
   DLY4X1 FE_PHC218_n1226 (.Y(FE_PHN218_n1226), 
	.A(FE_PHN5084_n1226));
   DLY4X1 FE_PHC217_n1295 (.Y(FE_PHN217_n1295), 
	.A(n1295));
   DLY4X1 FE_PHC216_n1260 (.Y(FE_PHN216_n1260), 
	.A(n1260));
   DLY4X1 FE_PHC215_n1323 (.Y(FE_PHN215_n1323), 
	.A(FE_PHN5123_n1323));
   DLY4X1 FE_PHC214_n1310 (.Y(FE_PHN214_n1310), 
	.A(n1310));
   DLY4X1 FE_PHC213_n1330 (.Y(FE_PHN213_n1330), 
	.A(n1330));
   DLY4X1 FE_PHC212_n1246 (.Y(FE_PHN212_n1246), 
	.A(n1246));
   DLY4X1 FE_PHC211_n1289 (.Y(FE_PHN211_n1289), 
	.A(FE_PHN5195_n1289));
   DLY4X1 FE_PHC210_n1314 (.Y(FE_PHN210_n1314), 
	.A(n1314));
   DLY4X1 FE_PHC209_n1250 (.Y(FE_PHN209_n1250), 
	.A(FE_PHN5175_n1250));
   DLY4X1 FE_PHC208_n1245 (.Y(FE_PHN208_n1245), 
	.A(FE_PHN5082_n1245));
   DLY4X1 FE_PHC207_n1247 (.Y(FE_PHN207_n1247), 
	.A(FE_PHN5186_n1247));
   DLY4X1 FE_PHC206_n1333 (.Y(FE_PHN206_n1333), 
	.A(n1333));
   DLY4X1 FE_PHC205_n1282 (.Y(FE_PHN205_n1282), 
	.A(n1282));
   DLY4X1 FE_PHC204_n1235 (.Y(FE_PHN204_n1235), 
	.A(n1235));
   DLY4X1 FE_PHC203_n1291 (.Y(FE_PHN203_n1291), 
	.A(FE_PHN5163_n1291));
   DLY4X1 FE_PHC202_n1325 (.Y(FE_PHN202_n1325), 
	.A(n1325));
   DLY4X1 FE_PHC201_n1219 (.Y(FE_PHN201_n1219), 
	.A(FE_PHN5166_n1219));
   DLY4X1 FE_PHC200_n1298 (.Y(FE_PHN200_n1298), 
	.A(n1298));
   DLY4X1 FE_PHC199_n1326 (.Y(FE_PHN199_n1326), 
	.A(FE_PHN5181_n1326));
   DLY4X1 FE_PHC197_n1320 (.Y(FE_PHN197_n1320), 
	.A(n1320));
   DLY4X1 FE_PHC196_n1279 (.Y(FE_PHN196_n1279), 
	.A(n1279));
   DLY4X1 FE_PHC195_n1278 (.Y(FE_PHN195_n1278), 
	.A(n1278));
   DLY4X1 FE_PHC194_n1256 (.Y(FE_PHN194_n1256), 
	.A(n1256));
   DLY4X1 FE_PHC193_n1263 (.Y(FE_PHN193_n1263), 
	.A(n1263));
   DLY4X1 FE_PHC192_n1294 (.Y(FE_PHN192_n1294), 
	.A(n1294));
   DLY4X1 FE_PHC191_n1293 (.Y(FE_PHN191_n1293), 
	.A(n1293));
   DLY4X1 FE_PHC190_n1242 (.Y(FE_PHN190_n1242), 
	.A(FE_PHN5182_n1242));
   DLY4X1 FE_PHC189_n1329 (.Y(FE_PHN189_n1329), 
	.A(n1329));
   DLY4X1 FE_PHC188_n1331 (.Y(FE_PHN188_n1331), 
	.A(n1331));
   DLY4X1 FE_PHC187_n1313 (.Y(FE_PHN187_n1313), 
	.A(n1313));
   DLY4X1 FE_PHC186_n1321 (.Y(FE_PHN186_n1321), 
	.A(n1321));
   DLY4X1 FE_PHC185_n1312 (.Y(FE_PHN185_n1312), 
	.A(n1312));
   DLY4X1 FE_PHC184_n1217 (.Y(FE_PHN184_n1217), 
	.A(n1217));
   DLY4X1 FE_PHC183_n1225 (.Y(FE_PHN183_n1225), 
	.A(n1225));
   DLY4X1 FE_PHC182_n1236 (.Y(FE_PHN182_n1236), 
	.A(FE_PHN5093_n1236));
   DLY4X1 FE_PHC181_n1266 (.Y(FE_PHN181_n1266), 
	.A(n1266));
   DLY4X1 FE_PHC180_n1230 (.Y(FE_PHN180_n1230), 
	.A(FE_PHN5120_n1230));
   DLY4X1 FE_PHC179_n1234 (.Y(FE_PHN179_n1234), 
	.A(FE_PHN5176_n1234));
   DLY4X1 FE_PHC177_n1220 (.Y(FE_PHN177_n1220), 
	.A(n1220));
   DLY4X1 FE_PHC176_n1315 (.Y(FE_PHN176_n1315), 
	.A(n1315));
   DLY4X1 FE_PHC175_n1283 (.Y(FE_PHN175_n1283), 
	.A(FE_PHN5222_n1283));
   DLY4X1 FE_PHC174_n1251 (.Y(FE_PHN174_n1251), 
	.A(n1251));
   DLY4X1 FE_PHC173_n1249 (.Y(FE_PHN173_n1249), 
	.A(FE_PHN5200_n1249));
   DLY4X1 FE_PHC172_n1218 (.Y(FE_PHN172_n1218), 
	.A(FE_PHN5188_n1218));
   DLY4X1 FE_PHC171_n1288 (.Y(FE_PHN171_n1288), 
	.A(n1288));
   DLY4X1 FE_PHC170_n1262 (.Y(FE_PHN170_n1262), 
	.A(n1262));
   DLY4X1 FE_PHC169_n1248 (.Y(FE_PHN169_n1248), 
	.A(FE_PHN5189_n1248));
   DLY4X1 FE_PHC168_n1261 (.Y(FE_PHN168_n1261), 
	.A(n1261));
   DLY4X1 FE_PHC167_n1299 (.Y(FE_PHN167_n1299), 
	.A(n1299));
   DLY4X1 FE_PHC166_n1328 (.Y(FE_PHN166_n1328), 
	.A(FE_PHN5194_n1328));
   DLY4X1 FE_PHC165_n1281 (.Y(FE_PHN165_n1281), 
	.A(FE_PHN5088_n1281));
   DLY4X1 FE_PHC164_n1233 (.Y(FE_PHN164_n1233), 
	.A(n1233));
   DLY4X1 FE_PHC163_n1280 (.Y(FE_PHN163_n1280), 
	.A(FE_PHN5190_n1280));
   DLY4X1 FE_PHC162_n1244 (.Y(FE_PHN162_n1244), 
	.A(FE_PHN5100_n1244));
   DLY4X1 FE_PHC161_n1297 (.Y(FE_PHN161_n1297), 
	.A(FE_PHN5169_n1297));
   DLY4X1 FE_PHC160_n1267 (.Y(FE_PHN160_n1267), 
	.A(FE_PHN5094_n1267));
   DLY4X1 FE_PHC159_n1265 (.Y(FE_PHN159_n1265), 
	.A(n1265));
   DLY4X1 FE_PHC158_n1264 (.Y(FE_PHN158_n1264), 
	.A(n1264));
   CLKBUFX3 FE_PHC157_n237 (.Y(FE_PHN157_n237), 
	.A(n237));
   DLY4X1 FE_PHC156_n1213 (.Y(FE_PHN156_n1213), 
	.A(FE_PHN5122_n1213));
   DLY4X1 FE_PHC154_n1308 (.Y(FE_PHN154_n1308), 
	.A(FE_PHN5118_n1308));
   DLY4X1 FE_PHC153_n1276 (.Y(FE_PHN153_n1276), 
	.A(FE_PHN5246_n1276));
   DLY4X1 FE_PHC152_n1237 (.Y(FE_PHN152_n1237), 
	.A(FE_PHN5135_n1237));
   DLY4X1 FE_PHC151_n1296 (.Y(FE_PHN151_n1296), 
	.A(FE_PHN5252_n1296));
   DLY4X1 FE_PHC150_n1257 (.Y(FE_PHN150_n1257), 
	.A(FE_PHN5191_n1257));
   DLY4X1 FE_PHC149_n1259 (.Y(FE_PHN149_n1259), 
	.A(n1259));
   DLY4X1 FE_PHC148_n1239 (.Y(FE_PHN148_n1239), 
	.A(FE_PHN5178_n1239));
   DLY4X1 FE_PHC147_n1207 (.Y(FE_PHN147_n1207), 
	.A(n1207));
   DLY4X1 FE_PHC146_n1206 (.Y(FE_PHN146_n1206), 
	.A(FE_PHN5140_n1206));
   DLY4X1 FE_PHC145_n1238 (.Y(FE_PHN145_n1238), 
	.A(FE_PHN5225_n1238));
   DLY4X1 FE_PHC144_n1269 (.Y(FE_PHN144_n1269), 
	.A(FE_PHN5179_n1269));
   DLY4X1 FE_PHC143_n1302 (.Y(FE_PHN143_n1302), 
	.A(n1302));
   DLY4X1 FE_PHC142_n1304 (.Y(FE_PHN142_n1304), 
	.A(FE_PHN5087_n1304));
   DLY4X1 FE_PHC141_n1301 (.Y(FE_PHN141_n1301), 
	.A(FE_PHN2806_n1301));
   DLY4X1 FE_PHC140_n1208 (.Y(FE_PHN140_n1208), 
	.A(FE_PHN5198_n1208));
   DLY4X1 FE_PHC139_n1303 (.Y(FE_PHN139_n1303), 
	.A(FE_PHN5115_n1303));
   DLY4X1 FE_PHC138_n1270 (.Y(FE_PHN138_n1270), 
	.A(n1270));
   DLY4X1 FE_PHC137_n1271 (.Y(FE_PHN137_n1271), 
	.A(n1271));
   DLY4X1 FE_PHC136_n1231 (.Y(FE_PHN136_n1231), 
	.A(n1231));
   DLY4X1 FE_PHC135_n1274 (.Y(FE_PHN135_n1274), 
	.A(FE_PHN5162_n1274));
   DLY4X1 FE_PHC134_n1211 (.Y(FE_PHN134_n1211), 
	.A(n1211));
   DLY4X1 FE_PHC133_n1241 (.Y(FE_PHN133_n1241), 
	.A(n1241));
   DLY4X1 FE_PHC132_n1243 (.Y(FE_PHN132_n1243), 
	.A(FE_PHN5099_n1243));
   DLY4X1 FE_PHC131_n1240 (.Y(FE_PHN131_n1240), 
	.A(FE_PHN5245_n1240));
   DLY4X1 FE_PHC130_n1209 (.Y(FE_PHN130_n1209), 
	.A(FE_PHN5203_n1209));
   DLY4X1 FE_PHC129_n1192 (.Y(FE_PHN129_n1192), 
	.A(n1192));
   DLY4X1 FE_PHC128_n1275 (.Y(FE_PHN128_n1275), 
	.A(n1275));
   DLY4X1 FE_PHC127_n1307 (.Y(FE_PHN127_n1307), 
	.A(FE_PHN5160_n1307));
   DLY4X1 FE_PHC126_n1210 (.Y(FE_PHN126_n1210), 
	.A(FE_PHN5130_n1210));
   DLY4X1 FE_PHC125_n1305 (.Y(FE_PHN125_n1305), 
	.A(n1305));
   DLY4X1 FE_PHC123_n1273 (.Y(FE_PHN123_n1273), 
	.A(FE_PHN5205_n1273));
   DLY4X1 FE_PHC122_n1306 (.Y(FE_PHN122_n1306), 
	.A(FE_PHN5090_n1306));
   DLY4X1 FE_PHC121_n1212 (.Y(FE_PHN121_n1212), 
	.A(FE_PHN5124_n1212));
   DLY4X1 FE_PHC118_n1272 (.Y(FE_PHN118_n1272), 
	.A(n1272));
   DLY4X1 FE_PHC117_n1268 (.Y(FE_PHN117_n1268), 
	.A(FE_PHN5247_n1268));
   DLY4X1 FE_PHC114_sword_ctr_reg_1_ (.Y(FE_PHN114_sword_ctr_reg_1_), 
	.A(sword_ctr_reg[1]));
   DLY4X1 FE_PHC113_n1189 (.Y(FE_PHN113_n1189), 
	.A(n1189));
   DLY4X1 FE_PHC111_enc_ctrl_reg_1_ (.Y(FE_PHN111_enc_ctrl_reg_1_), 
	.A(enc_ctrl_reg[1]));
   CLKBUFX2 FE_OFC98_n232 (.Y(FE_OFN98_n232), 
	.A(FE_OFN97_n232));
   CLKBUFX3 FE_OFC97_n232 (.Y(FE_OFN97_n232), 
	.A(n232));
   DFFSX1 ready_reg_reg (.SN(FE_OFN39_reset_n), 
	.QN(), 
	.Q(ready), 
	.D(FE_PHN1310_n1334), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 block_w0_reg_reg_15_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN528_Dout_111_), 
	.D(FE_PHN249_n1222), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w0_reg_reg_23_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN3095_Dout_119_), 
	.D(FE_PHN226_n1214), 
	.CK(clk_48Mhz__L6_N44));
   JKFFRXL round_ctr_reg_reg_0_ (.RN(FE_OFN55_reset_n), 
	.QN(n54), 
	.Q(round[0]), 
	.K(n1201), 
	.J(FE_PHN3408_enc_ctrl_reg_0_), 
	.CK(clk));
   DFFRHQX1 block_w2_reg_reg_15_ (.RN(reset_n), 
	.Q(FE_PHN3105_Dout_47_), 
	.D(FE_PHN235_n1285), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w0_reg_reg_31_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN361_Dout_127_), 
	.D(FE_PHN146_n1206), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 block_w0_reg_reg_7_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN750_Dout_103_), 
	.D(FE_PHN180_n1230), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w3_reg_reg_15_ (.RN(reset_n), 
	.Q(FE_PHN336_Dout_15_), 
	.D(FE_PHN246_n1317), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w3_reg_reg_23_ (.RN(reset_n), 
	.Q(FE_PHN299_Dout_23_), 
	.D(FE_PHN221_n1309), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w2_reg_reg_23_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN300_Dout_55_), 
	.D(FE_PHN225_n1277), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w3_reg_reg_31_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN281_Dout_31_), 
	.D(FE_PHN141_n1301), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 block_w2_reg_reg_31_ (.RN(reset_n), 
	.Q(FE_PHN414_Dout_63_), 
	.D(FE_PHN144_n1269), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w2_reg_reg_7_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN378_Dout_39_), 
	.D(FE_PHN191_n1293), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w1_reg_reg_15_ (.RN(reset_n), 
	.Q(FE_PHN341_Dout_79_), 
	.D(FE_PHN233_n1253), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w1_reg_reg_23_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN278_Dout_87_), 
	.D(FE_PHN208_n1245), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w1_reg_reg_31_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN304_Dout_95_), 
	.D(FE_PHN152_n1237), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w1_reg_reg_7_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN269_Dout_71_), 
	.D(FE_PHN168_n1261), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 block_w0_reg_reg_14_ (.RN(reset_n), 
	.Q(FE_PHN595_Dout_110_), 
	.D(FE_PHN250_n1223), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w2_reg_reg_6_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN702_Dout_38_), 
	.D(FE_PHN192_n1294), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w2_reg_reg_14_ (.RN(reset_n), 
	.Q(FE_PHN601_Dout_46_), 
	.D(FE_PHN232_n1286), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 block_w0_reg_reg_30_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN412_Dout_126_), 
	.D(FE_PHN147_n1207), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 block_w3_reg_reg_14_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN295_Dout_14_), 
	.D(FE_PHN242_n1318), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 block_w2_reg_reg_22_ (.RN(reset_n), 
	.Q(FE_PHN440_Dout_54_), 
	.D(FE_PHN195_n1278), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w1_reg_reg_6_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN309_Dout_70_), 
	.D(FE_PHN170_n1262), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w1_reg_reg_14_ (.RN(reset_n), 
	.Q(FE_PHN292_Dout_78_), 
	.D(FE_PHN237_n1254), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w3_reg_reg_30_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN282_Dout_30_), 
	.D(FE_PHN5145_n1302), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 block_w2_reg_reg_30_ (.RN(reset_n), 
	.Q(FE_PHN318_Dout_62_), 
	.D(FE_PHN5196_n1270), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 block_w1_reg_reg_30_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN288_Dout_94_), 
	.D(FE_PHN145_n1238), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w1_reg_reg_22_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN279_Dout_86_), 
	.D(FE_PHN212_n1246), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w3_reg_reg_7_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN298_Dout_7_), 
	.D(FE_PHN202_n1325), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 block_w0_reg_reg_6_ (.RN(reset_n), 
	.Q(FE_PHN599_Dout_102_), 
	.D(FE_PHN136_n1231), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w3_reg_reg_6_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN377_Dout_6_), 
	.D(FE_PHN199_n1326), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 block_w0_reg_reg_22_ (.RN(reset_n), 
	.Q(FE_PHN330_Dout_118_), 
	.D(FE_PHN222_n1215), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 block_w3_reg_reg_22_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN365_Dout_22_), 
	.D(FE_PHN214_n1310), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 block_w2_reg_reg_2_ (.RN(FE_OFN56_reset_n), 
	.Q(FE_PHN604_Dout_34_), 
	.D(FE_PHN200_n1298), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 block_w0_reg_reg_26_ (.RN(FE_OFN55_reset_n), 
	.Q(FE_PHN533_Dout_122_), 
	.D(FE_PHN5095_n1211), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 block_w1_reg_reg_2_ (.RN(FE_OFN56_reset_n), 
	.Q(FE_PHN273_Dout_66_), 
	.D(FE_PHN5217_n1266), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w1_reg_reg_10_ (.RN(FE_OFN56_reset_n), 
	.Q(FE_PHN368_Dout_74_), 
	.D(FE_PHN227_n1258), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w1_reg_reg_11_ (.RN(reset_n), 
	.Q(FE_PHN293_Dout_75_), 
	.D(FE_PHN150_n1257), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w2_reg_reg_10_ (.RN(FE_OFN56_reset_n), 
	.Q(FE_PHN315_Dout_42_), 
	.D(FE_PHN5081_n1290), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w2_reg_reg_18_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN312_Dout_50_), 
	.D(FE_PHN5183_n1282), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w3_reg_reg_26_ (.RN(FE_OFN55_reset_n), 
	.Q(FE_PHN356_Dout_26_), 
	.D(FE_PHN122_n1306), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 block_w1_reg_reg_29_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN415_Dout_93_), 
	.D(FE_PHN148_n1239), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w1_reg_reg_18_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN274_Dout_82_), 
	.D(FE_PHN209_n1250), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w2_reg_reg_26_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN355_Dout_58_), 
	.D(FE_PHN135_n1274), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w1_reg_reg_26_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN321_Dout_90_), 
	.D(FE_PHN190_n1242), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w0_reg_reg_13_ (.RN(reset_n), 
	.Q(FE_PHN435_Dout_109_), 
	.D(FE_PHN243_n1224), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 block_w0_reg_reg_1_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN3106_Dout_97_), 
	.D(FE_PHN5248_n1236), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w0_reg_reg_5_ (.RN(reset_n), 
	.Q(FE_PHN596_Dout_101_), 
	.D(FE_PHN219_n1232), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 block_w3_reg_reg_1_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN821_Dout_1_), 
	.D(FE_PHN5249_n1331), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w3_reg_reg_8_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN3104_Dout_8_), 
	.D(FE_PHN5177_n1324), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w3_reg_reg_0_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN438_Dout_0_), 
	.D(FE_PHN247_n1332), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w0_reg_reg_10_ (.RN(FE_OFN55_reset_n), 
	.Q(new_block[106]), 
	.D(FE_PHN231_n1227), 
	.CK(clk));
   DFFRHQX1 block_w3_reg_reg_3_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN363_Dout_3_), 
	.D(FE_PHN5215_n1329), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w3_reg_reg_2_ (.RN(FE_OFN55_reset_n), 
	.Q(new_block[2]), 
	.D(FE_PHN2807_n1330), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w3_reg_reg_10_ (.RN(FE_OFN56_reset_n), 
	.Q(FE_PHN603_Dout_10_), 
	.D(FE_PHN244_n1322), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w2_reg_reg_5_ (.RN(reset_n), 
	.Q(FE_PHN600_Dout_37_), 
	.D(FE_PHN217_n1295), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w2_reg_reg_4_ (.RN(reset_n), 
	.Q(FE_PHN701_Dout_36_), 
	.D(FE_PHN151_n1296), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w2_reg_reg_13_ (.RN(reset_n), 
	.Q(FE_PHN362_Dout_45_), 
	.D(FE_PHN240_n1287), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w2_reg_reg_12_ (.RN(reset_n), 
	.Q(FE_PHN597_Dout_44_), 
	.D(FE_PHN171_n1288), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w2_reg_reg_1_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN3107_Dout_33_), 
	.D(FE_PHN5079_n1299), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w0_reg_reg_29_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN2850_Dout_125_), 
	.D(FE_PHN140_n1208), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 block_w3_reg_reg_5_ (.RN(reset_n), 
	.Q(FE_PHN259_Dout_5_), 
	.D(FE_PHN224_n1327), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 block_w3_reg_reg_13_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN307_Dout_13_), 
	.D(FE_PHN238_n1319), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 block_w0_reg_reg_21_ (.RN(reset_n), 
	.Q(FE_PHN436_Dout_117_), 
	.D(FE_PHN229_n1216), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 block_w0_reg_reg_3_ (.RN(reset_n), 
	.Q(FE_PHN311_Dout_99_), 
	.D(FE_PHN179_n1234), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w0_reg_reg_2_ (.RN(FE_OFN55_reset_n), 
	.Q(FE_PHN266_Dout_98_), 
	.D(FE_PHN5185_n1235), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w3_reg_reg_21_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN364_Dout_21_), 
	.D(FE_PHN220_n1311), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 block_w0_reg_reg_17_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN328_Dout_113_), 
	.D(FE_PHN5107_n1220), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w3_reg_reg_17_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN331_Dout_17_), 
	.D(FE_PHN5106_n1315), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w0_reg_reg_11_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN339_Dout_107_), 
	.D(FE_PHN218_n1226), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w3_reg_reg_11_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN338_Dout_11_), 
	.D(FE_PHN186_n1321), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w2_reg_reg_3_ (.RN(reset_n), 
	.Q(FE_PHN371_Dout_35_), 
	.D(FE_PHN161_n1297), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w2_reg_reg_0_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN313_Dout_32_), 
	.D(FE_PHN228_n1300), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w0_reg_reg_24_ (.RN(FE_OFN55_reset_n), 
	.Q(FE_PHN413_Dout_120_), 
	.D(FE_PHN156_n1213), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 block_w0_reg_reg_25_ (.RN(FE_OFN55_reset_n), 
	.Q(FE_PHN351_Dout_121_), 
	.D(FE_PHN121_n1212), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 block_w3_reg_reg_19_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN317_Dout_19_), 
	.D(FE_PHN187_n1313), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w3_reg_reg_16_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN310_Dout_16_), 
	.D(FE_PHN248_n1316), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w0_reg_reg_18_ (.RN(FE_OFN55_reset_n), 
	.Q(FE_PHN442_Dout_114_), 
	.D(FE_PHN201_n1219), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 block_w3_reg_reg_18_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN314_Dout_18_), 
	.D(FE_PHN5121_n1314), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w2_reg_reg_9_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN305_Dout_41_), 
	.D(FE_PHN203_n1291), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w2_reg_reg_21_ (.RN(reset_n), 
	.Q(FE_PHN374_Dout_53_), 
	.D(FE_PHN5218_n1279), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w2_reg_reg_17_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN334_Dout_49_), 
	.D(FE_PHN175_n1283), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w1_reg_reg_1_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN340_Dout_65_), 
	.D(FE_PHN160_n1267), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w1_reg_reg_4_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN373_Dout_68_), 
	.D(FE_PHN5250_n1264), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w1_reg_reg_5_ (.RN(reset_n), 
	.Q(FE_PHN261_Dout_69_), 
	.D(FE_PHN193_n1263), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w1_reg_reg_0_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN297_Dout_64_), 
	.D(FE_PHN117_n1268), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 block_w1_reg_reg_12_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN367_Dout_76_), 
	.D(FE_PHN5253_n1256), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w1_reg_reg_8_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN443_Dout_72_), 
	.D(FE_PHN216_n1260), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 block_w1_reg_reg_3_ (.RN(reset_n), 
	.Q(FE_PHN276_Dout_67_), 
	.D(FE_PHN5192_n1265), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w1_reg_reg_13_ (.RN(reset_n), 
	.Q(FE_PHN294_Dout_77_), 
	.D(FE_PHN234_n1255), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 block_w1_reg_reg_9_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN444_Dout_73_), 
	.D(FE_PHN149_n1259), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 block_w3_reg_reg_29_ (.RN(reset_n), 
	.Q(FE_PHN257_Dout_29_), 
	.D(FE_PHN139_n1303), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 block_w0_reg_reg_27_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN352_Dout_123_), 
	.D(FE_PHN126_n1210), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w2_reg_reg_11_ (.RN(reset_n), 
	.Q(FE_PHN260_Dout_43_), 
	.D(FE_PHN211_n1289), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w2_reg_reg_19_ (.RN(reset_n), 
	.Q(FE_PHN306_Dout_51_), 
	.D(FE_PHN165_n1281), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w2_reg_reg_8_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN280_Dout_40_), 
	.D(FE_PHN236_n1292), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w2_reg_reg_16_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN333_Dout_48_), 
	.D(FE_PHN239_n1284), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w3_reg_reg_24_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN286_Dout_24_), 
	.D(FE_PHN154_n1308), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 block_w3_reg_reg_25_ (.RN(FE_OFN55_reset_n), 
	.Q(FE_PHN285_Dout_25_), 
	.D(FE_PHN127_n1307), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 block_w2_reg_reg_28_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN353_Dout_60_), 
	.D(FE_PHN5202_n1272), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w2_reg_reg_29_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN262_Dout_61_), 
	.D(FE_PHN137_n1271), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 block_w2_reg_reg_25_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN284_Dout_57_), 
	.D(FE_PHN5111_n1275), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w1_reg_reg_28_ (.RN(reset_n), 
	.Q(FE_PHN303_Dout_92_), 
	.D(FE_PHN131_n1240), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w1_reg_reg_19_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN267_Dout_83_), 
	.D(FE_PHN173_n1249), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w1_reg_reg_21_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN316_Dout_85_), 
	.D(FE_PHN207_n1247), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w1_reg_reg_16_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN308_Dout_80_), 
	.D(FE_PHN5219_n1252), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w1_reg_reg_17_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN277_Dout_81_), 
	.D(FE_PHN5136_n1251), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w3_reg_reg_27_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN264_Dout_27_), 
	.D(FE_PHN5143_n1305), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 block_w2_reg_reg_24_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN263_Dout_56_), 
	.D(FE_PHN153_n1276), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w2_reg_reg_27_ (.RN(reset_n), 
	.Q(FE_PHN287_Dout_59_), 
	.D(FE_PHN123_n1273), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w1_reg_reg_24_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN320_Dout_88_), 
	.D(FE_PHN5216_n1244), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w1_reg_reg_25_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN272_Dout_89_), 
	.D(FE_PHN132_n1243), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w1_reg_reg_27_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN289_Dout_91_), 
	.D(FE_PHN5226_n1241), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w0_reg_reg_4_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN433_Dout_100_), 
	.D(FE_PHN5187_n1233), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w0_reg_reg_12_ (.RN(reset_n), 
	.Q(FE_PHN437_Dout_108_), 
	.D(FE_PHN5201_n1225), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w0_reg_reg_8_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN3108_Dout_104_), 
	.D(FE_PHN251_n1229), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w0_reg_reg_9_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN369_Dout_105_), 
	.D(FE_PHN223_n1228), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w3_reg_reg_4_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN329_Dout_4_), 
	.D(FE_PHN166_n1328), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w3_reg_reg_9_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN441_Dout_9_), 
	.D(FE_PHN215_n1323), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 block_w0_reg_reg_20_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN598_Dout_116_), 
	.D(FE_PHN184_n1217), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w3_reg_reg_20_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN366_Dout_20_), 
	.D(FE_PHN185_n1312), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w0_reg_reg_28_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN350_Dout_124_), 
	.D(FE_PHN130_n1209), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w0_reg_reg_0_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN268_Dout_96_), 
	.D(FE_PHN5097_n1333), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 block_w3_reg_reg_12_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN275_Dout_12_), 
	.D(FE_PHN197_n1320), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w0_reg_reg_16_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN335_Dout_112_), 
	.D(FE_PHN5096_n1221), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 block_w0_reg_reg_19_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN337_Dout_115_), 
	.D(FE_PHN172_n1218), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w2_reg_reg_20_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN332_Dout_52_), 
	.D(FE_PHN163_n1280), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w3_reg_reg_28_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN302_Dout_28_), 
	.D(FE_PHN142_n1304), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 block_w1_reg_reg_20_ (.RN(FE_OFN54_reset_n), 
	.Q(FE_PHN296_Dout_84_), 
	.D(FE_PHN169_n1248), 
	.CK(clk_48Mhz__L6_N41));
   JKFFRXL sword_ctr_reg_reg_0_ (.RN(FE_OFN55_reset_n), 
	.QN(n56), 
	.Q(sword_ctr_reg[0]), 
	.K(n1203), 
	.J(n1193), 
	.CK(clk));
   DFFRHQX1 sword_ctr_reg_reg_1_ (.RN(FE_OFN55_reset_n), 
	.Q(sword_ctr_reg[1]), 
	.D(FE_PHN2809_n1340), 
	.CK(clk));
   DFFRHQX1 enc_ctrl_reg_reg_1_ (.RN(FE_OFN55_reset_n), 
	.Q(enc_ctrl_reg[1]), 
	.D(FE_PHN258_n1339), 
	.CK(clk));
   DFFRHQX1 enc_ctrl_reg_reg_0_ (.RN(FE_OFN39_reset_n), 
	.Q(enc_ctrl_reg[0]), 
	.D(FE_PHN2856_n1338), 
	.CK(clk));
   DFFRHQX1 round_ctr_reg_reg_3_ (.RN(FE_OFN55_reset_n), 
	.Q(round[3]), 
	.D(FE_PHN354_n1335), 
	.CK(clk));
   DFFRHQX1 round_ctr_reg_reg_1_ (.RN(FE_OFN55_reset_n), 
	.Q(FE_PHN2812_enc_round_nr_1_), 
	.D(FE_PHN751_n1337), 
	.CK(clk));
   DFFRHQX1 round_ctr_reg_reg_2_ (.RN(FE_OFN39_reset_n), 
	.Q(round[2]), 
	.D(FE_PHN703_n1336), 
	.CK(clk));
   NAND2X1 U3 (.Y(n1), 
	.B(n230), 
	.A(n702));
   NAND2X1 U4 (.Y(n2), 
	.B(n706), 
	.A(n702));
   NAND2X1 U5 (.Y(n3), 
	.B(n945), 
	.A(n702));
   INVX1 U8 (.Y(n30), 
	.A(n35));
   INVX2 U10 (.Y(n105), 
	.A(n111));
   INVX2 U15 (.Y(n9), 
	.A(n228));
   INVX1 U16 (.Y(n15), 
	.A(n227));
   NOR3X1 U18 (.Y(n703), 
	.C(n93), 
	.B(n110), 
	.A(FE_OFN98_n232));
   INVX1 U21 (.Y(n13), 
	.A(n1));
   INVX1 U22 (.Y(n12), 
	.A(n1));
   INVX1 U23 (.Y(n17), 
	.A(n2));
   INVX1 U24 (.Y(n8), 
	.A(n3));
   INVX1 U25 (.Y(n7), 
	.A(n3));
   INVX1 U26 (.Y(n16), 
	.A(n2));
   INVX1 U27 (.Y(n11), 
	.A(n464));
   INVX2 U31 (.Y(n106), 
	.A(n110));
   INVX2 U32 (.Y(n107), 
	.A(n110));
   INVX1 U39 (.Y(n108), 
	.A(n110));
   INVX1 U41 (.Y(n111), 
	.A(n99));
   INVX1 U43 (.Y(n113), 
	.A(n105));
   INVX1 U44 (.Y(n114), 
	.A(n107));
   INVX1 U47 (.Y(n35), 
	.A(FE_PHN157_n237));
   INVX1 U52 (.Y(n48), 
	.A(FE_PHN157_n237));
   INVX1 U60 (.Y(n47), 
	.A(FE_PHN157_n237));
   INVX1 U63 (.Y(n51), 
	.A(FE_PHN157_n237));
   INVX1 U67 (.Y(n49), 
	.A(FE_PHN157_n237));
   INVX1 U69 (.Y(n50), 
	.A(FE_PHN157_n237));
   INVX1 U71 (.Y(n46), 
	.A(FE_PHN157_n237));
   INVX1 U83 (.Y(n38), 
	.A(FE_PHN157_n237));
   INVX1 U86 (.Y(n39), 
	.A(FE_PHN157_n237));
   INVX1 U92 (.Y(n14), 
	.A(n227));
   NAND2X2 U93 (.Y(n945), 
	.B(n193), 
	.A(n703));
   INVX1 U104 (.Y(n93), 
	.A(FE_PHN157_n237));
   INVX1 U105 (.Y(n110), 
	.A(n236));
   INVX1 U107 (.Y(n99), 
	.A(n110));
   INVX1 U110 (.Y(n83), 
	.A(FE_PHN157_n237));
   INVX1 U122 (.Y(n173), 
	.A(n228));
   INVX1 U126 (.Y(n141), 
	.A(new_sboxw[26]));
   INVX1 U127 (.Y(n138), 
	.A(new_sboxw[29]));
   INVX1 U128 (.Y(n139), 
	.A(new_sboxw[31]));
   INVX1 U129 (.Y(n137), 
	.A(new_sboxw[30]));
   INVX1 U130 (.Y(n143), 
	.A(new_sboxw[24]));
   INVX1 U131 (.Y(n142), 
	.A(new_sboxw[25]));
   INVX1 U132 (.Y(n140), 
	.A(new_sboxw[28]));
   INVX1 U133 (.Y(n144), 
	.A(new_sboxw[27]));
   NOR2X1 U134 (.Y(n232), 
	.B(n1190), 
	.A(n176));
   NAND2X2 U135 (.Y(n706), 
	.B(n227), 
	.A(n703));
   NAND2X2 U136 (.Y(n465), 
	.B(n228), 
	.A(n703));
   NAND2X2 U137 (.Y(n230), 
	.B(n194), 
	.A(n703));
   AND2X2 U138 (.Y(n4), 
	.B(n465), 
	.A(n702));
   INVX1 U139 (.Y(n464), 
	.A(n4));
   INVX2 U144 (.Y(n97), 
	.A(FE_PHN157_n237));
   CLKINVX3 U145 (.Y(n96), 
	.A(FE_PHN157_n237));
   NOR2X1 U146 (.Y(n702), 
	.B(n1190), 
	.A(FE_PHN113_n1189));
   AOI21X1 U147 (.Y(n1191), 
	.B0(n183), 
	.A1(n181), 
	.A0(n182));
   AOI2BB1X1 U148 (.Y(n1190), 
	.B0(n1193), 
	.A1N(FE_PHN129_n1192), 
	.A0N(n1191));
   NAND2X1 U149 (.Y(n227), 
	.B(n702), 
	.A(FE_PHN256_n943));
   NAND2X1 U150 (.Y(n228), 
	.B(n702), 
	.A(FE_PHN253_n704));
   NAND2X2 U151 (.Y(n193), 
	.B(n702), 
	.A(n1182));
   NAND2X1 U154 (.Y(n236), 
	.B(FE_PHN113_n1189), 
	.A(n1190));
   INVX1 U155 (.Y(n176), 
	.A(FE_PHN113_n1189));
   INVX1 U156 (.Y(n151), 
	.A(round_key[59]));
   INVX1 U157 (.Y(n150), 
	.A(round_key[91]));
   INVX1 U158 (.Y(n152), 
	.A(round_key[27]));
   INVX1 U159 (.Y(n149), 
	.A(round_key[123]));
   INVX1 U160 (.Y(n148), 
	.A(round_key[26]));
   INVX1 U161 (.Y(n145), 
	.A(round_key[122]));
   INVX1 U162 (.Y(n146), 
	.A(round_key[90]));
   INVX1 U163 (.Y(n147), 
	.A(round_key[58]));
   INVX1 U164 (.Y(n135), 
	.A(round_key[57]));
   INVX1 U165 (.Y(n136), 
	.A(round_key[25]));
   INVX1 U166 (.Y(n133), 
	.A(round_key[121]));
   INVX1 U167 (.Y(n134), 
	.A(round_key[89]));
   INVX1 U168 (.Y(n166), 
	.A(round_key[88]));
   INVX1 U169 (.Y(n168), 
	.A(round_key[24]));
   INVX1 U170 (.Y(n165), 
	.A(round_key[120]));
   INVX1 U171 (.Y(n169), 
	.A(round_key[127]));
   INVX1 U172 (.Y(n162), 
	.A(round_key[94]));
   INVX1 U173 (.Y(n161), 
	.A(round_key[126]));
   INVX1 U174 (.Y(n157), 
	.A(round_key[125]));
   INVX1 U175 (.Y(n158), 
	.A(round_key[93]));
   INVX1 U176 (.Y(n154), 
	.A(round_key[92]));
   INVX1 U177 (.Y(n167), 
	.A(round_key[56]));
   INVX1 U178 (.Y(n171), 
	.A(round_key[63]));
   INVX1 U179 (.Y(n163), 
	.A(round_key[62]));
   INVX1 U180 (.Y(n159), 
	.A(round_key[61]));
   INVX1 U181 (.Y(n155), 
	.A(round_key[60]));
   INVX1 U182 (.Y(n156), 
	.A(round_key[28]));
   INVX1 U183 (.Y(n153), 
	.A(round_key[124]));
   INVX1 U184 (.Y(n172), 
	.A(round_key[31]));
   INVX1 U185 (.Y(n164), 
	.A(round_key[30]));
   INVX1 U186 (.Y(n160), 
	.A(round_key[29]));
   INVX1 U187 (.Y(n170), 
	.A(round_key[95]));
   NAND2BX4 U189 (.Y(n237), 
	.B(n1191), 
	.AN(FE_PHN129_n1192));
   XNOR2X1 U190 (.Y(n936), 
	.B(n1359), 
	.A(round_key[33]));
   XNOR2X1 U191 (.Y(n1160), 
	.B(n1396), 
	.A(round_key[3]));
   XNOR2X1 U192 (.Y(n338), 
	.B(n1441), 
	.A(round_key[115]));
   XNOR2X1 U193 (.Y(n1065), 
	.B(n1369), 
	.A(round_key[17]));
   XNOR2X1 U194 (.Y(n353), 
	.B(n1427), 
	.A(round_key[113]));
   XNOR2X1 U195 (.Y(n585), 
	.B(n1425), 
	.A(round_key[81]));
   XNOR2X1 U196 (.Y(n826), 
	.B(n1437), 
	.A(round_key[49]));
   XNOR2X1 U197 (.Y(n803), 
	.B(n1388), 
	.A(round_key[52]));
   XNOR2X1 U198 (.Y(n1050), 
	.B(n1371), 
	.A(round_key[19]));
   XNOR2X1 U199 (.Y(n1175), 
	.B(n1434), 
	.A(round_key[1]));
   XNOR2X1 U200 (.Y(n1042), 
	.B(n1396), 
	.A(round_key[20]));
   XNOR2X1 U201 (.Y(n330), 
	.B(n1383), 
	.A(round_key[116]));
   XNOR2X1 U202 (.Y(n570), 
	.B(n1449), 
	.A(round_key[83]));
   XNOR2X1 U203 (.Y(n448), 
	.B(n1345), 
	.A(round_key[99]));
   XNOR2X1 U204 (.Y(n680), 
	.B(n1395), 
	.A(round_key[67]));
   XNOR2X1 U205 (.Y(n440), 
	.B(n1374), 
	.A(round_key[100]));
   XNOR2X1 U206 (.Y(n562), 
	.B(n1399), 
	.A(round_key[84]));
   XNOR2X1 U207 (.Y(n811), 
	.B(n1450), 
	.A(round_key[51]));
   XNOR2X1 U208 (.Y(n672), 
	.B(n1382), 
	.A(round_key[68]));
   XNOR2X1 U209 (.Y(n913), 
	.B(n1373), 
	.A(round_key[36]));
   XNOR2X1 U210 (.Y(n463), 
	.B(n1360), 
	.A(round_key[97]));
   XNOR2X1 U211 (.Y(n1152), 
	.B(n1365), 
	.A(round_key[4]));
   XNOR2X1 U212 (.Y(n921), 
	.B(n1344), 
	.A(round_key[35]));
   XNOR2X1 U213 (.Y(n695), 
	.B(n1370), 
	.A(round_key[65]));
   XOR2X1 U214 (.Y(n1164), 
	.B(n1166), 
	.A(n1165));
   XNOR2X1 U215 (.Y(n1166), 
	.B(n987), 
	.A(n1435));
   XNOR2X1 U216 (.Y(n1165), 
	.B(n1167), 
	.A(n1453));
   XNOR2X1 U217 (.Y(n1167), 
	.B(n1371), 
	.A(round_key[2]));
   XOR2X1 U218 (.Y(n925), 
	.B(n927), 
	.A(n926));
   XNOR2X1 U219 (.Y(n927), 
	.B(n748), 
	.A(n1361));
   XNOR2X1 U220 (.Y(n926), 
	.B(n928), 
	.A(n1437));
   XNOR2X1 U221 (.Y(n928), 
	.B(n185), 
	.A(round_key[34]));
   XOR2X1 U222 (.Y(n1054), 
	.B(n1056), 
	.A(n1055));
   XNOR2X1 U223 (.Y(n1056), 
	.B(n995), 
	.A(n1432));
   XNOR2X1 U224 (.Y(n1055), 
	.B(n1057), 
	.A(n1444));
   XNOR2X1 U225 (.Y(n1057), 
	.B(n1434), 
	.A(round_key[18]));
   XOR2X1 U226 (.Y(n574), 
	.B(n576), 
	.A(n575));
   XNOR2X1 U227 (.Y(n576), 
	.B(n515), 
	.A(n1428));
   XNOR2X1 U228 (.Y(n575), 
	.B(n577), 
	.A(n1440));
   XNOR2X1 U229 (.Y(n577), 
	.B(n1370), 
	.A(round_key[82]));
   XOR2X1 U230 (.Y(n1016), 
	.B(n1018), 
	.A(n1017));
   XNOR2X1 U231 (.Y(n1018), 
	.B(n1019), 
	.A(n1407));
   XNOR2X1 U232 (.Y(n1017), 
	.B(n1020), 
	.A(n1367));
   XNOR2X1 U233 (.Y(n1020), 
	.B(n1379), 
	.A(round_key[23]));
   XOR2X1 U234 (.Y(n647), 
	.B(n649), 
	.A(n648));
   XNOR2X1 U235 (.Y(n649), 
	.B(n473), 
	.A(n1354));
   XNOR2X1 U236 (.Y(n648), 
	.B(n650), 
	.A(n1410));
   XNOR2X1 U237 (.Y(n650), 
	.B(n1358), 
	.A(round_key[71]));
   XOR2X1 U238 (.Y(n684), 
	.B(n686), 
	.A(n685));
   XNOR2X1 U239 (.Y(n686), 
	.B(n507), 
	.A(n1455));
   XNOR2X1 U240 (.Y(n685), 
	.B(n687), 
	.A(n1429));
   XNOR2X1 U241 (.Y(n687), 
	.B(n1343), 
	.A(round_key[66]));
   XOR2X1 U242 (.Y(n888), 
	.B(n890), 
	.A(n889));
   XNOR2X1 U243 (.Y(n890), 
	.B(n714), 
	.A(n1390));
   XNOR2X1 U244 (.Y(n889), 
	.B(n891), 
	.A(n1391));
   XNOR2X1 U245 (.Y(n891), 
	.B(n1355), 
	.A(round_key[39]));
   XOR2X1 U246 (.Y(n634), 
	.B(n636), 
	.A(n635));
   XOR2X1 U247 (.Y(n636), 
	.B(n616), 
	.A(n532));
   XOR2X1 U248 (.Y(n635), 
	.B(n637), 
	.A(n516));
   XNOR2X1 U249 (.Y(n637), 
	.B(n1343), 
	.A(round_key[73]));
   XOR2X1 U250 (.Y(n1114), 
	.B(n1116), 
	.A(n1115));
   XOR2X1 U251 (.Y(n1116), 
	.B(n1096), 
	.A(n1012));
   XOR2X1 U252 (.Y(n1115), 
	.B(n1117), 
	.A(n996));
   XNOR2X1 U253 (.Y(n1117), 
	.B(n1453), 
	.A(round_key[9]));
   XOR2X1 U254 (.Y(n875), 
	.B(n877), 
	.A(n876));
   XOR2X1 U255 (.Y(n877), 
	.B(n857), 
	.A(n773));
   XOR2X1 U256 (.Y(n876), 
	.B(n878), 
	.A(n757));
   XNOR2X1 U257 (.Y(n878), 
	.B(n185), 
	.A(round_key[41]));
   XOR2X1 U258 (.Y(n1108), 
	.B(n1110), 
	.A(n1109));
   XOR2X1 U259 (.Y(n1110), 
	.B(n1003), 
	.A(n987));
   XNOR2X1 U260 (.Y(n1109), 
	.B(n1451), 
	.A(round_key[10]));
   XOR2X1 U261 (.Y(n589), 
	.B(n591), 
	.A(n590));
   XOR2X1 U262 (.Y(n591), 
	.B(n532), 
	.A(n473));
   XNOR2X1 U263 (.Y(n590), 
	.B(n1426), 
	.A(round_key[80]));
   XOR2X1 U264 (.Y(n1121), 
	.B(n1123), 
	.A(n1122));
   XOR2X1 U265 (.Y(n1123), 
	.B(n1096), 
	.A(n1004));
   XNOR2X1 U266 (.Y(n1122), 
	.B(n1393), 
	.A(round_key[8]));
   XOR2X1 U267 (.Y(n830), 
	.B(n832), 
	.A(n831));
   XOR2X1 U268 (.Y(n832), 
	.B(n773), 
	.A(n714));
   XNOR2X1 U269 (.Y(n831), 
	.B(n1392), 
	.A(round_key[48]));
   XOR2X1 U270 (.Y(n1069), 
	.B(n1071), 
	.A(n1070));
   XOR2X1 U271 (.Y(n1071), 
	.B(n1012), 
	.A(n953));
   XNOR2X1 U272 (.Y(n1070), 
	.B(n1422), 
	.A(round_key[16]));
   XOR2X1 U273 (.Y(n882), 
	.B(n884), 
	.A(n883));
   XOR2X1 U274 (.Y(n884), 
	.B(n857), 
	.A(n765));
   XNOR2X1 U275 (.Y(n883), 
	.B(n1359), 
	.A(round_key[40]));
   XOR2X1 U276 (.Y(n409), 
	.B(n411), 
	.A(n410));
   XOR2X1 U277 (.Y(n411), 
	.B(n384), 
	.A(n292));
   XNOR2X1 U278 (.Y(n410), 
	.B(n1342), 
	.A(round_key[104]));
   XOR2X1 U279 (.Y(n940), 
	.B(n942), 
	.A(n941));
   XOR2X1 U280 (.Y(n942), 
	.B(n780), 
	.A(n765));
   XNOR2X1 U281 (.Y(n941), 
	.B(n1419), 
	.A(round_key[32]));
   XOR2X1 U282 (.Y(n641), 
	.B(n643), 
	.A(n642));
   XOR2X1 U283 (.Y(n643), 
	.B(n616), 
	.A(n524));
   XNOR2X1 U284 (.Y(n642), 
	.B(n184), 
	.A(round_key[72]));
   XOR2X1 U285 (.Y(n396), 
	.B(n398), 
	.A(n397));
   XOR2X1 U286 (.Y(n398), 
	.B(n291), 
	.A(n275));
   XNOR2X1 U287 (.Y(n397), 
	.B(n1454), 
	.A(round_key[106]));
   XOR2X1 U288 (.Y(n1179), 
	.B(n1181), 
	.A(n1180));
   XOR2X1 U289 (.Y(n1181), 
	.B(n1019), 
	.A(n1004));
   XNOR2X1 U290 (.Y(n1180), 
	.B(n1369), 
	.A(round_key[0]));
   XOR2X1 U291 (.Y(n375), 
	.B(n377), 
	.A(n376));
   XOR2X1 U292 (.Y(n377), 
	.B(n266), 
	.A(n249));
   XNOR2X1 U293 (.Y(n376), 
	.B(n192), 
	.A(round_key[109]));
   XOR2X1 U294 (.Y(n621), 
	.B(n623), 
	.A(n622));
   XOR2X1 U295 (.Y(n623), 
	.B(n616), 
	.A(n515));
   XOR2X1 U296 (.Y(n622), 
	.B(n624), 
	.A(n496));
   XNOR2X1 U297 (.Y(n624), 
	.B(n1382), 
	.A(round_key[75]));
   XOR2X1 U298 (.Y(n1101), 
	.B(n1103), 
	.A(n1102));
   XOR2X1 U299 (.Y(n1103), 
	.B(n1096), 
	.A(n995));
   XOR2X1 U300 (.Y(n1102), 
	.B(n1104), 
	.A(n976));
   XNOR2X1 U301 (.Y(n1104), 
	.B(n188), 
	.A(round_key[11]));
   XOR2X1 U302 (.Y(n862), 
	.B(n864), 
	.A(n863));
   XOR2X1 U303 (.Y(n864), 
	.B(n857), 
	.A(n756));
   XOR2X1 U304 (.Y(n863), 
	.B(n865), 
	.A(n737));
   XNOR2X1 U305 (.Y(n865), 
	.B(n1373), 
	.A(round_key[43]));
   XNOR2X1 U306 (.Y(n1178), 
	.B(n1393), 
	.A(round_key[0]));
   XOR2X1 U307 (.Y(n357), 
	.B(n359), 
	.A(n358));
   XOR2X1 U308 (.Y(n359), 
	.B(n300), 
	.A(n241));
   XNOR2X1 U309 (.Y(n358), 
	.B(n1418), 
	.A(round_key[112]));
   XOR2X1 U310 (.Y(n342), 
	.B(n344), 
	.A(n343));
   XNOR2X1 U311 (.Y(n344), 
	.B(n283), 
	.A(n1442));
   XNOR2X1 U312 (.Y(n343), 
	.B(n345), 
	.A(n1360));
   XNOR2X1 U313 (.Y(n345), 
	.B(n1430), 
	.A(round_key[114]));
   XOR2X1 U314 (.Y(n815), 
	.B(n817), 
	.A(n816));
   XNOR2X1 U315 (.Y(n817), 
	.B(n756), 
	.A(n1433));
   XNOR2X1 U316 (.Y(n816), 
	.B(n818), 
	.A(n1436));
   XNOR2X1 U317 (.Y(n818), 
	.B(n1438), 
	.A(round_key[50]));
   XOR2X1 U318 (.Y(n402), 
	.B(n404), 
	.A(n403));
   XOR2X1 U319 (.Y(n404), 
	.B(n384), 
	.A(n300));
   XOR2X1 U320 (.Y(n403), 
	.B(n405), 
	.A(n284));
   XNOR2X1 U321 (.Y(n405), 
	.B(n1394), 
	.A(round_key[105]));
   XOR2X1 U322 (.Y(n304), 
	.B(n306), 
	.A(n305));
   XNOR2X1 U323 (.Y(n306), 
	.B(n307), 
	.A(n1353));
   XNOR2X1 U324 (.Y(n305), 
	.B(n308), 
	.A(n1356));
   XNOR2X1 U325 (.Y(n308), 
	.B(n1411), 
	.A(round_key[119]));
   XOR2X1 U326 (.Y(n536), 
	.B(n538), 
	.A(n537));
   XNOR2X1 U327 (.Y(n538), 
	.B(n539), 
	.A(n1378));
   XNOR2X1 U328 (.Y(n537), 
	.B(n540), 
	.A(n1368));
   XNOR2X1 U329 (.Y(n540), 
	.B(n1409), 
	.A(round_key[87]));
   XOR2X1 U330 (.Y(n777), 
	.B(n779), 
	.A(n778));
   XNOR2X1 U331 (.Y(n779), 
	.B(n780), 
	.A(n229));
   XNOR2X1 U332 (.Y(n778), 
	.B(n781), 
	.A(n1199));
   XNOR2X1 U333 (.Y(n781), 
	.B(n1408), 
	.A(round_key[55]));
   XOR2X1 U334 (.Y(n544), 
	.B(n546), 
	.A(n545));
   XNOR2X1 U335 (.Y(n546), 
	.B(n480), 
	.A(n1366));
   XNOR2X1 U336 (.Y(n545), 
	.B(n547), 
	.A(n1403));
   XNOR2X1 U337 (.Y(n547), 
	.B(n1410), 
	.A(round_key[86]));
   XOR2X1 U338 (.Y(n785), 
	.B(n787), 
	.A(n786));
   XNOR2X1 U339 (.Y(n787), 
	.B(n721), 
	.A(n190));
   XNOR2X1 U340 (.Y(n786), 
	.B(n788), 
	.A(n1402));
   XNOR2X1 U341 (.Y(n788), 
	.B(n1390), 
	.A(round_key[54]));
   XOR2X1 U342 (.Y(n1024), 
	.B(n1026), 
	.A(n1025));
   XNOR2X1 U343 (.Y(n1026), 
	.B(n960), 
	.A(n1375));
   XNOR2X1 U344 (.Y(n1025), 
	.B(n1027), 
	.A(n1377));
   XNOR2X1 U345 (.Y(n1027), 
	.B(n1401), 
	.A(round_key[22]));
   XOR2X1 U346 (.Y(n312), 
	.B(n314), 
	.A(n313));
   XNOR2X1 U347 (.Y(n314), 
	.B(n248), 
	.A(n1406));
   XNOR2X1 U348 (.Y(n313), 
	.B(n315), 
	.A(n1350));
   XNOR2X1 U349 (.Y(n315), 
	.B(n1404), 
	.A(round_key[118]));
   XOR2X1 U350 (.Y(n551), 
	.B(n553), 
	.A(n552));
   XNOR2X1 U351 (.Y(n553), 
	.B(n488), 
	.A(n1348));
   XNOR2X1 U352 (.Y(n552), 
	.B(n554), 
	.A(n1398));
   XNOR2X1 U353 (.Y(n554), 
	.B(n1400), 
	.A(round_key[85]));
   XOR2X1 U354 (.Y(n792), 
	.B(n794), 
	.A(n793));
   XNOR2X1 U355 (.Y(n794), 
	.B(n729), 
	.A(n1346));
   XNOR2X1 U356 (.Y(n793), 
	.B(n795), 
	.A(n1387));
   XNOR2X1 U357 (.Y(n795), 
	.B(n1389), 
	.A(round_key[53]));
   XOR2X1 U358 (.Y(n1031), 
	.B(n1033), 
	.A(n1032));
   XNOR2X1 U359 (.Y(n1033), 
	.B(n968), 
	.A(n1385));
   XNOR2X1 U360 (.Y(n1032), 
	.B(n1034), 
	.A(n1376));
   XNOR2X1 U361 (.Y(n1034), 
	.B(n1365), 
	.A(round_key[21]));
   XOR2X1 U362 (.Y(n607), 
	.B(n609), 
	.A(n608));
   XOR2X1 U363 (.Y(n609), 
	.B(n498), 
	.A(n481));
   XNOR2X1 U364 (.Y(n608), 
	.B(n1351), 
	.A(round_key[77]));
   XOR2X1 U365 (.Y(n452), 
	.B(n454), 
	.A(n453));
   XNOR2X1 U366 (.Y(n454), 
	.B(n275), 
	.A(n1431));
   XNOR2X1 U367 (.Y(n453), 
	.B(n455), 
	.A(n1394));
   XNOR2X1 U368 (.Y(n455), 
	.B(n186), 
	.A(round_key[98]));
   XOR2X1 U369 (.Y(n1127), 
	.B(n1129), 
	.A(n1128));
   XNOR2X1 U370 (.Y(n1129), 
	.B(n953), 
	.A(n1377));
   XNOR2X1 U371 (.Y(n1128), 
	.B(n1130), 
	.A(n1380));
   XNOR2X1 U372 (.Y(n1130), 
	.B(n705), 
	.A(round_key[7]));
   XOR2X1 U373 (.Y(n595), 
	.B(n597), 
	.A(n596));
   XOR2X1 U374 (.Y(n597), 
	.B(n539), 
	.A(n480));
   XNOR2X1 U375 (.Y(n596), 
	.B(n1413), 
	.A(round_key[79]));
   XOR2X1 U376 (.Y(n1081), 
	.B(n1083), 
	.A(n1082));
   XOR2X1 U377 (.Y(n1083), 
	.B(n968), 
	.A(n952));
   XNOR2X1 U378 (.Y(n1082), 
	.B(n705), 
	.A(round_key[14]));
   XOR2X1 U379 (.Y(n319), 
	.B(n321), 
	.A(n320));
   XNOR2X1 U380 (.Y(n321), 
	.B(n256), 
	.A(n1405));
   XNOR2X1 U381 (.Y(n320), 
	.B(n322), 
	.A(n1374));
   XNOR2X1 U382 (.Y(n322), 
	.B(n1363), 
	.A(round_key[117]));
   XOR2X1 U383 (.Y(n854), 
	.B(n856), 
	.A(n855));
   XOR2X1 U384 (.Y(n856), 
	.B(n857), 
	.A(n747));
   XOR2X1 U385 (.Y(n855), 
	.B(n858), 
	.A(n730));
   XNOR2X1 U386 (.Y(n858), 
	.B(n1349), 
	.A(round_key[44]));
   XOR2X1 U387 (.Y(n628), 
	.B(n630), 
	.A(n629));
   XOR2X1 U388 (.Y(n630), 
	.B(n523), 
	.A(n507));
   XNOR2X1 U389 (.Y(n629), 
	.B(n1395), 
	.A(round_key[74]));
   XOR2X1 U390 (.Y(n1075), 
	.B(n1077), 
	.A(n1076));
   XOR2X1 U391 (.Y(n1077), 
	.B(n1019), 
	.A(n960));
   XNOR2X1 U392 (.Y(n1076), 
	.B(n1415), 
	.A(round_key[15]));
   XOR2X1 U393 (.Y(n601), 
	.B(n603), 
	.A(n602));
   XOR2X1 U394 (.Y(n603), 
	.B(n488), 
	.A(n472));
   XNOR2X1 U395 (.Y(n602), 
	.B(n1354), 
	.A(round_key[78]));
   XOR2X1 U396 (.Y(n1087), 
	.B(n1089), 
	.A(n1088));
   XOR2X1 U397 (.Y(n1089), 
	.B(n978), 
	.A(n961));
   XNOR2X1 U398 (.Y(n1088), 
	.B(n191), 
	.A(round_key[13]));
   XOR2X1 U399 (.Y(n613), 
	.B(n615), 
	.A(n614));
   XOR2X1 U400 (.Y(n615), 
	.B(n616), 
	.A(n506));
   XOR2X1 U401 (.Y(n614), 
	.B(n617), 
	.A(n489));
   XNOR2X1 U402 (.Y(n617), 
	.B(n1364), 
	.A(round_key[76]));
   XOR2X1 U403 (.Y(n699), 
	.B(n701), 
	.A(n700));
   XOR2X1 U404 (.Y(n701), 
	.B(n539), 
	.A(n524));
   XNOR2X1 U405 (.Y(n700), 
	.B(n1425), 
	.A(round_key[64]));
   XOR2X1 U406 (.Y(n415), 
	.B(n417), 
	.A(n416));
   XNOR2X1 U407 (.Y(n417), 
	.B(n241), 
	.A(n1406));
   XNOR2X1 U408 (.Y(n416), 
	.B(n418), 
	.A(n1417));
   XNOR2X1 U409 (.Y(n418), 
	.B(n944), 
	.A(round_key[103]));
   XOR2X1 U410 (.Y(n836), 
	.B(n838), 
	.A(n837));
   XOR2X1 U411 (.Y(n838), 
	.B(n780), 
	.A(n721));
   XNOR2X1 U412 (.Y(n837), 
	.B(n1416), 
	.A(round_key[47]));
   XOR2X1 U413 (.Y(n654), 
	.B(n656), 
	.A(n655));
   XNOR2X1 U414 (.Y(n656), 
	.B(n472), 
	.A(n1351));
   XNOR2X1 U415 (.Y(n655), 
	.B(n657), 
	.A(n1378));
   XNOR2X1 U416 (.Y(n657), 
	.B(n1400), 
	.A(round_key[70]));
   XOR2X1 U417 (.Y(n422), 
	.B(n424), 
	.A(n423));
   XNOR2X1 U418 (.Y(n424), 
	.B(n240), 
	.A(n1405));
   XNOR2X1 U419 (.Y(n423), 
	.B(n425), 
	.A(n1353));
   XNOR2X1 U420 (.Y(n425), 
	.B(n192), 
	.A(round_key[102]));
   XOR2X1 U421 (.Y(n842), 
	.B(n844), 
	.A(n843));
   XOR2X1 U422 (.Y(n844), 
	.B(n729), 
	.A(n713));
   XNOR2X1 U423 (.Y(n843), 
	.B(n1355), 
	.A(round_key[46]));
   XOR2X1 U424 (.Y(n661), 
	.B(n663), 
	.A(n662));
   XNOR2X1 U425 (.Y(n663), 
	.B(n481), 
	.A(n1364));
   XNOR2X1 U426 (.Y(n662), 
	.B(n664), 
	.A(n1366));
   XNOR2X1 U427 (.Y(n664), 
	.B(n1399), 
	.A(round_key[69]));
   XOR2X1 U428 (.Y(n429), 
	.B(n431), 
	.A(n430));
   XNOR2X1 U429 (.Y(n431), 
	.B(n249), 
	.A(n1384));
   XNOR2X1 U430 (.Y(n430), 
	.B(n432), 
	.A(n1350));
   XNOR2X1 U431 (.Y(n432), 
	.B(n189), 
	.A(round_key[101]));
   XOR2X1 U432 (.Y(n848), 
	.B(n850), 
	.A(n849));
   XOR2X1 U433 (.Y(n850), 
	.B(n739), 
	.A(n722));
   XNOR2X1 U434 (.Y(n849), 
	.B(n1352), 
	.A(round_key[45]));
   XOR2X1 U435 (.Y(n1093), 
	.B(n1095), 
	.A(n1094));
   XOR2X1 U436 (.Y(n1095), 
	.B(n1096), 
	.A(n986));
   XOR2X1 U437 (.Y(n1094), 
	.B(n1097), 
	.A(n969));
   XNOR2X1 U438 (.Y(n1097), 
	.B(n1347), 
	.A(round_key[12]));
   XOR2X1 U439 (.Y(n381), 
	.B(n383), 
	.A(n382));
   XOR2X1 U440 (.Y(n383), 
	.B(n384), 
	.A(n274));
   XOR2X1 U441 (.Y(n382), 
	.B(n385), 
	.A(n257));
   XNOR2X1 U442 (.Y(n385), 
	.B(n189), 
	.A(round_key[108]));
   XOR2X1 U443 (.Y(n363), 
	.B(n365), 
	.A(n364));
   XOR2X1 U444 (.Y(n365), 
	.B(n307), 
	.A(n248));
   XNOR2X1 U445 (.Y(n364), 
	.B(n1414), 
	.A(round_key[111]));
   XOR2X1 U446 (.Y(n1134), 
	.B(n1136), 
	.A(n1135));
   XNOR2X1 U447 (.Y(n1136), 
	.B(n952), 
	.A(n1376));
   XNOR2X1 U448 (.Y(n1135), 
	.B(n1137), 
	.A(n191));
   XNOR2X1 U449 (.Y(n1137), 
	.B(n1367), 
	.A(round_key[6]));
   XOR2X1 U450 (.Y(n895), 
	.B(n897), 
	.A(n896));
   XNOR2X1 U451 (.Y(n897), 
	.B(n713), 
	.A(n229));
   XNOR2X1 U452 (.Y(n896), 
	.B(n898), 
	.A(n1389));
   XNOR2X1 U453 (.Y(n898), 
	.B(n1352), 
	.A(round_key[38]));
   XOR2X1 U454 (.Y(n369), 
	.B(n371), 
	.A(n370));
   XOR2X1 U455 (.Y(n371), 
	.B(n256), 
	.A(n240));
   XNOR2X1 U456 (.Y(n370), 
	.B(n944), 
	.A(round_key[110]));
   XOR2X1 U457 (.Y(n1141), 
	.B(n1143), 
	.A(n1142));
   XNOR2X1 U458 (.Y(n1143), 
	.B(n961), 
	.A(n1386));
   XNOR2X1 U459 (.Y(n1142), 
	.B(n1144), 
	.A(n1347));
   XNOR2X1 U460 (.Y(n1144), 
	.B(n1401), 
	.A(round_key[5]));
   XOR2X1 U461 (.Y(n902), 
	.B(n904), 
	.A(n903));
   XNOR2X1 U462 (.Y(n904), 
	.B(n722), 
	.A(n190));
   XNOR2X1 U463 (.Y(n903), 
	.B(n905), 
	.A(n1388));
   XNOR2X1 U464 (.Y(n905), 
	.B(n1349), 
	.A(round_key[37]));
   XOR2X1 U465 (.Y(n389), 
	.B(n391), 
	.A(n390));
   XOR2X1 U466 (.Y(n391), 
	.B(n384), 
	.A(n283));
   XOR2X1 U467 (.Y(n390), 
	.B(n392), 
	.A(n264));
   XNOR2X1 U468 (.Y(n392), 
	.B(n1452), 
	.A(round_key[107]));
   XOR2X1 U469 (.Y(n869), 
	.B(n871), 
	.A(n870));
   XOR2X1 U470 (.Y(n871), 
	.B(n764), 
	.A(n748));
   XNOR2X1 U471 (.Y(n870), 
	.B(n1344), 
	.A(round_key[42]));
   XOR2X1 U472 (.Y(n1186), 
	.B(n1188), 
	.A(n1187));
   XOR2X1 U473 (.Y(n1188), 
	.B(n307), 
	.A(n292));
   XNOR2X1 U474 (.Y(n1187), 
	.B(n1420), 
	.A(round_key[96]));
   NAND2X1 U475 (.Y(n1201), 
	.B(FE_PHN3081_n1194), 
	.A(n180));
   INVX1 U476 (.Y(n179), 
	.A(FE_PHN602_n1197));
   OAI211X1 U477 (.Y(n1338), 
	.C0(n1202), 
	.B0(FE_PHN3081_n1194), 
	.A1(n180), 
	.A0(FE_PHN535_enc_ctrl_we));
   OAI211X1 U478 (.Y(n1339), 
	.C0(n1202), 
	.B0(n176), 
	.A1(n178), 
	.A0(FE_PHN535_enc_ctrl_we));
   NAND2X1 U479 (.Y(n1203), 
	.B(n177), 
	.A(n180));
   INVX1 U480 (.Y(n177), 
	.A(n1193));
   NAND2X1 U481 (.Y(n1202), 
	.B(FE_PHN535_enc_ctrl_we), 
	.A(n1193));
   OAI21XL U482 (.Y(n1340), 
	.B0(n1204), 
	.A1(n1203), 
	.A0(n175));
   OAI21XL U483 (.Y(n1204), 
	.B0(n1193), 
	.A1(FE_PHN256_n943), 
	.A0(FE_PHN253_n704));
   OAI22X1 U484 (.Y(n1189), 
	.B1(FE_PHN129_n1192), 
	.B0(n1191), 
	.A1(n180), 
	.A0(FE_PHN111_enc_ctrl_reg_1_));
   INVX1 U485 (.Y(n181), 
	.A(round[1]));
   INVX1 U486 (.Y(n182), 
	.A(FE_PHN2813_enc_round_nr_2_));
   INVX1 U487 (.Y(n183), 
	.A(round[3]));
   NAND3X2 U488 (.Y(n194), 
	.C(n702), 
	.B(n175), 
	.A(n56));
   AOI22X1 U489 (.Y(n206), 
	.B1(n15), 
	.B0(new_block[60]), 
	.A1(n9), 
	.A0(new_block[92]));
   AOI22X1 U490 (.Y(n214), 
	.B1(n15), 
	.B0(new_block[52]), 
	.A1(n9), 
	.A0(FE_PHN296_Dout_84_));
   AOI22X1 U491 (.Y(n200), 
	.B1(n15), 
	.B0(FE_PHN701_Dout_36_), 
	.A1(n9), 
	.A0(new_block[68]));
   OAI221XL U492 (.Y(sboxw[28]), 
	.C0(n206), 
	.B1(n1384), 
	.B0(n194), 
	.A1(n1386), 
	.A0(n193));
   OAI221XL U493 (.Y(sboxw[20]), 
	.C0(n214), 
	.B1(n1385), 
	.B0(n194), 
	.A1(n1387), 
	.A0(n193));
   OAI221XL U494 (.Y(sboxw[4]), 
	.C0(n200), 
	.B1(n1364), 
	.B0(n194), 
	.A1(n189), 
	.A0(n193));
   INVX1 U495 (.Y(n180), 
	.A(FE_PHN3408_enc_ctrl_reg_0_));
   NOR2X1 U496 (.Y(n1193), 
	.B(n178), 
	.A(FE_PHN3408_enc_ctrl_reg_0_));
   OAI221XL U497 (.Y(sboxw[24]), 
	.C0(n210), 
	.B1(n1418), 
	.B0(n194), 
	.A1(n1422), 
	.A0(n193));
   AOI22X1 U498 (.Y(n210), 
	.B1(n15), 
	.B0(new_block[56]), 
	.A1(n9), 
	.A0(new_block[88]));
   INVX1 U499 (.Y(n178), 
	.A(FE_PHN2821_enc_ctrl_reg_1_));
   NAND2X1 U500 (.Y(n1192), 
	.B(FE_PHN111_enc_ctrl_reg_1_), 
	.A(FE_PHN3408_enc_ctrl_reg_0_));
   AOI22X1 U501 (.Y(n207), 
	.B1(n15), 
	.B0(new_block[59]), 
	.A1(n9), 
	.A0(new_block[91]));
   AOI22X1 U502 (.Y(n205), 
	.B1(n15), 
	.B0(new_block[61]), 
	.A1(n9), 
	.A0(new_block[93]));
   AOI22X1 U503 (.Y(n224), 
	.B1(n14), 
	.B0(FE_PHN260_Dout_43_), 
	.A1(n173), 
	.A0(FE_PHN293_Dout_75_));
   AOI22X1 U504 (.Y(n216), 
	.B1(n14), 
	.B0(new_block[51]), 
	.A1(n9), 
	.A0(new_block[83]));
   AOI22X1 U505 (.Y(n217), 
	.B1(n14), 
	.B0(new_block[50]), 
	.A1(n173), 
	.A0(new_block[82]));
   AOI22X1 U506 (.Y(n196), 
	.B1(n15), 
	.B0(new_block[40]), 
	.A1(n9), 
	.A0(new_block[72]));
   AOI22X1 U507 (.Y(n225), 
	.B1(n14), 
	.B0(FE_PHN315_Dout_42_), 
	.A1(n173), 
	.A0(new_block[74]));
   OAI221XL U508 (.Y(sboxw[8]), 
	.C0(n196), 
	.B1(n1419), 
	.B0(n194), 
	.A1(n1425), 
	.A0(n193));
   AOI22X1 U509 (.Y(n213), 
	.B1(n15), 
	.B0(new_block[53]), 
	.A1(n9), 
	.A0(FE_PHN316_Dout_85_));
   OAI221XL U510 (.Y(sboxw[10]), 
	.C0(n225), 
	.B1(n1361), 
	.B0(n194), 
	.A1(n1455), 
	.A0(n193));
   OAI221XL U511 (.Y(sboxw[18]), 
	.C0(n217), 
	.B1(n1443), 
	.B0(n194), 
	.A1(n1445), 
	.A0(n193));
   OAI221XL U512 (.Y(sboxw[2]), 
	.C0(n204), 
	.B1(n1395), 
	.B0(n194), 
	.A1(n1454), 
	.A0(n193));
   AOI22X1 U513 (.Y(n195), 
	.B1(n15), 
	.B0(FE_PHN305_Dout_41_), 
	.A1(n9), 
	.A0(new_block[73]));
   AOI22X1 U514 (.Y(n222), 
	.B1(n14), 
	.B0(FE_PHN362_Dout_45_), 
	.A1(n173), 
	.A0(FE_PHN294_Dout_77_));
   AOI22X1 U515 (.Y(n204), 
	.B1(n15), 
	.B0(new_block[34]), 
	.A1(n9), 
	.A0(new_block[66]));
   AOI22X1 U516 (.Y(n223), 
	.B1(n14), 
	.B0(FE_PHN597_Dout_44_), 
	.A1(n173), 
	.A0(FE_PHN367_Dout_76_));
   AOI22X1 U517 (.Y(n199), 
	.B1(n15), 
	.B0(FE_PHN600_Dout_37_), 
	.A1(n9), 
	.A0(new_block[69]));
   AOI22X1 U518 (.Y(n201), 
	.B1(n15), 
	.B0(FE_PHN371_Dout_35_), 
	.A1(n9), 
	.A0(new_block[67]));
   OAI221XL U519 (.Y(sboxw[12]), 
	.C0(n223), 
	.B1(n1346), 
	.B0(n194), 
	.A1(n1348), 
	.A0(n193));
   OAI221XL U520 (.Y(sboxw[25]), 
	.C0(n209), 
	.B1(n1431), 
	.B0(n194), 
	.A1(n1435), 
	.A0(n193));
   AOI22X1 U521 (.Y(n209), 
	.B1(n15), 
	.B0(new_block[57]), 
	.A1(n9), 
	.A0(new_block[89]));
   OAI221XL U522 (.Y(sboxw[16]), 
	.C0(n219), 
	.B1(n1421), 
	.B0(n194), 
	.A1(n1423), 
	.A0(n193));
   AOI22X1 U523 (.Y(n219), 
	.B1(n14), 
	.B0(new_block[48]), 
	.A1(n173), 
	.A0(FE_PHN308_Dout_80_));
   OAI221XL U524 (.Y(sboxw[0]), 
	.C0(n226), 
	.B1(n184), 
	.B0(n194), 
	.A1(n1342), 
	.A0(n193));
   AOI22X1 U525 (.Y(n226), 
	.B1(n14), 
	.B0(new_block[32]), 
	.A1(n173), 
	.A0(new_block[64]));
   OAI221XL U526 (.Y(sboxw[17]), 
	.C0(n218), 
	.B1(n1432), 
	.B0(n194), 
	.A1(n1436), 
	.A0(n193));
   AOI22X1 U527 (.Y(n218), 
	.B1(n14), 
	.B0(new_block[49]), 
	.A1(n173), 
	.A0(FE_PHN277_Dout_81_));
   OAI221XL U528 (.Y(sboxw[1]), 
	.C0(n215), 
	.B1(n1343), 
	.B0(n194), 
	.A1(n1394), 
	.A0(n193));
   AOI22X1 U529 (.Y(n215), 
	.B1(n14), 
	.B0(new_block[33]), 
	.A1(n173), 
	.A0(new_block[65]));
   OAI221XL U530 (.Y(sboxw[9]), 
	.C0(n195), 
	.B1(n1433), 
	.B0(n194), 
	.A1(n1370), 
	.A0(n193));
   OAI221XL U531 (.Y(sboxw[11]), 
	.C0(n224), 
	.B1(n187), 
	.B0(n194), 
	.A1(n1372), 
	.A0(n193));
   OAI221XL U532 (.Y(sboxw[27]), 
	.C0(n207), 
	.B1(n1446), 
	.B0(n194), 
	.A1(n1448), 
	.A0(n193));
   OAI221XL U533 (.Y(sboxw[19]), 
	.C0(n216), 
	.B1(n1447), 
	.B0(n194), 
	.A1(n1397), 
	.A0(n193));
   OAI221XL U534 (.Y(sboxw[3]), 
	.C0(n201), 
	.B1(n1382), 
	.B0(n194), 
	.A1(n1452), 
	.A0(n193));
   OAI221XL U535 (.Y(sboxw[5]), 
	.C0(n199), 
	.B1(n1351), 
	.B0(n194), 
	.A1(n192), 
	.A0(n193));
   OAI221XL U536 (.Y(sboxw[13]), 
	.C0(n222), 
	.B1(n190), 
	.B0(n194), 
	.A1(n1366), 
	.A0(n193));
   OAI221XL U537 (.Y(sboxw[29]), 
	.C0(n205), 
	.B1(n1405), 
	.B0(n194), 
	.A1(n1376), 
	.A0(n193));
   OAI221XL U538 (.Y(sboxw[21]), 
	.C0(n213), 
	.B1(n1375), 
	.B0(n194), 
	.A1(n1402), 
	.A0(n193));
   OAI221XL U539 (.Y(n1322), 
	.C0(n1106), 
	.B1(n945), 
	.B0(n1455), 
	.A1(n108), 
	.A0(n1105));
   XNOR2X1 U540 (.Y(n1105), 
	.B(block[10]), 
	.A(round_key[10]));
   AOI222X1 U541 (.Y(n1106), 
	.C1(n1108), 
	.C0(FE_OFN98_n232), 
	.B1(n1107), 
	.B0(n96), 
	.A1(new_sboxw[10]), 
	.A0(n7));
   XNOR2X1 U542 (.Y(n1107), 
	.B(n1371), 
	.A(round_key[10]));
   OAI221XL U543 (.Y(n1330), 
	.C0(n1162), 
	.B1(n945), 
	.B0(n1454), 
	.A1(n108), 
	.A0(n1161));
   XNOR2X1 U544 (.Y(n1161), 
	.B(block[2]), 
	.A(round_key[2]));
   AOI222X1 U545 (.Y(n1162), 
	.C1(n1164), 
	.C0(n232), 
	.B1(n1163), 
	.B0(n96), 
	.A1(new_sboxw[2]), 
	.A0(n7));
   XNOR2X1 U546 (.Y(n1163), 
	.B(n1451), 
	.A(round_key[2]));
   OAI221XL U547 (.Y(n1298), 
	.C0(n923), 
	.B1(n706), 
	.B0(n1451), 
	.A1(n107), 
	.A0(n922));
   XNOR2X1 U548 (.Y(n922), 
	.B(block[34]), 
	.A(round_key[34]));
   AOI222X1 U549 (.Y(n923), 
	.C1(n925), 
	.C0(FE_OFN98_n232), 
	.B1(n924), 
	.B0(n97), 
	.A1(new_sboxw[2]), 
	.A0(n16));
   XNOR2X1 U550 (.Y(n924), 
	.B(n1344), 
	.A(round_key[34]));
   OAI221XL U551 (.Y(n1314), 
	.C0(n1052), 
	.B1(n945), 
	.B0(n1445), 
	.A1(n107), 
	.A0(n1051));
   XNOR2X1 U552 (.Y(n1051), 
	.B(block[18]), 
	.A(round_key[18]));
   AOI222X1 U553 (.Y(n1052), 
	.C1(n1054), 
	.C0(n232), 
	.B1(n1053), 
	.B0(n83), 
	.A1(new_sboxw[18]), 
	.A0(n8));
   XNOR2X1 U554 (.Y(n1053), 
	.B(n1443), 
	.A(round_key[18]));
   OAI221XL U555 (.Y(n1250), 
	.C0(n572), 
	.B1(n465), 
	.B0(n1441), 
	.A1(n106), 
	.A0(n571));
   XNOR2X1 U556 (.Y(n571), 
	.B(block[82]), 
	.A(round_key[82]));
   AOI222X1 U557 (.Y(n572), 
	.C1(n574), 
	.C0(FE_OFN98_n232), 
	.B1(n573), 
	.B0(n47), 
	.A1(new_sboxw[18]), 
	.A0(n11));
   XNOR2X1 U558 (.Y(n573), 
	.B(n1439), 
	.A(round_key[82]));
   OAI221XL U559 (.Y(n1282), 
	.C0(n813), 
	.B1(n706), 
	.B0(n1439), 
	.A1(n106), 
	.A0(n812));
   XNOR2X1 U560 (.Y(n812), 
	.B(block[50]), 
	.A(round_key[50]));
   AOI222X1 U561 (.Y(n813), 
	.C1(n815), 
	.C0(FE_OFN98_n232), 
	.B1(n814), 
	.B0(n83), 
	.A1(new_sboxw[18]), 
	.A0(n17));
   XNOR2X1 U562 (.Y(n814), 
	.B(n1445), 
	.A(round_key[50]));
   OAI221XL U563 (.Y(n1309), 
	.C0(n1014), 
	.B1(n945), 
	.B0(n1416), 
	.A1(n107), 
	.A0(FE_PHN2816_n1013));
   XNOR2X1 U564 (.Y(n1013), 
	.B(block[23]), 
	.A(round_key[23]));
   AOI222X1 U565 (.Y(n1014), 
	.C1(n1016), 
	.C0(FE_OFN97_n232), 
	.B1(n1015), 
	.B0(n97), 
	.A1(new_sboxw[23]), 
	.A0(n8));
   XNOR2X1 U566 (.Y(n1015), 
	.B(n1415), 
	.A(round_key[23]));
   OAI221XL U567 (.Y(n1245), 
	.C0(n534), 
	.B1(n465), 
	.B0(n1414), 
	.A1(n99), 
	.A0(n533));
   XNOR2X1 U568 (.Y(n533), 
	.B(block[87]), 
	.A(round_key[87]));
   AOI222X1 U569 (.Y(n534), 
	.C1(n536), 
	.C0(FE_OFN97_n232), 
	.B1(n535), 
	.B0(n96), 
	.A1(new_sboxw[23]), 
	.A0(n11));
   XNOR2X1 U570 (.Y(n535), 
	.B(n1413), 
	.A(round_key[87]));
   OAI221XL U571 (.Y(n1277), 
	.C0(n775), 
	.B1(n706), 
	.B0(n1413), 
	.A1(n236), 
	.A0(FE_PHN5214_n774));
   XNOR2X1 U572 (.Y(n774), 
	.B(block[55]), 
	.A(round_key[55]));
   AOI222X1 U573 (.Y(n775), 
	.C1(n777), 
	.C0(FE_OFN97_n232), 
	.B1(n776), 
	.B0(n96), 
	.A1(new_sboxw[23]), 
	.A0(n17));
   XNOR2X1 U574 (.Y(n776), 
	.B(n1416), 
	.A(round_key[55]));
   OAI221XL U575 (.Y(n1261), 
	.C0(n645), 
	.B1(n465), 
	.B0(n1412), 
	.A1(n236), 
	.A0(n644));
   XNOR2X1 U576 (.Y(n644), 
	.B(block[71]), 
	.A(round_key[71]));
   AOI222X1 U577 (.Y(n645), 
	.C1(n647), 
	.C0(FE_OFN97_n232), 
	.B1(n646), 
	.B0(n96), 
	.A1(new_sboxw[7]), 
	.A0(n4));
   XNOR2X1 U578 (.Y(n646), 
	.B(n1357), 
	.A(round_key[71]));
   OAI221XL U579 (.Y(n1325), 
	.C0(n1125), 
	.B1(n945), 
	.B0(n1381), 
	.A1(n108), 
	.A0(n1124));
   XNOR2X1 U580 (.Y(n1124), 
	.B(block[7]), 
	.A(round_key[7]));
   AOI222X1 U581 (.Y(n1125), 
	.C1(n1127), 
	.C0(FE_OFN97_n232), 
	.B1(n1126), 
	.B0(n96), 
	.A1(new_sboxw[7]), 
	.A0(n7));
   XNOR2X1 U582 (.Y(n1126), 
	.B(n1341), 
	.A(round_key[7]));
   OAI221XL U583 (.Y(n1258), 
	.C0(n626), 
	.B1(n465), 
	.B0(n1371), 
	.A1(n106), 
	.A0(n625));
   XNOR2X1 U584 (.Y(n625), 
	.B(block[74]), 
	.A(round_key[74]));
   AOI222X1 U585 (.Y(n626), 
	.C1(n628), 
	.C0(FE_OFN98_n232), 
	.B1(n627), 
	.B0(n51), 
	.A1(new_sboxw[10]), 
	.A0(n4));
   XNOR2X1 U586 (.Y(n627), 
	.B(n1455), 
	.A(round_key[74]));
   OAI221XL U587 (.Y(n1263), 
	.C0(n659), 
	.B1(n465), 
	.B0(n1352), 
	.A1(n236), 
	.A0(FE_PHN5235_n658));
   XNOR2X1 U588 (.Y(n658), 
	.B(block[69]), 
	.A(round_key[69]));
   AOI222X1 U589 (.Y(n659), 
	.C1(n661), 
	.C0(FE_OFN97_n232), 
	.B1(n660), 
	.B0(n96), 
	.A1(new_sboxw[5]), 
	.A0(n4));
   XNOR2X1 U590 (.Y(n660), 
	.B(n1351), 
	.A(round_key[69]));
   OAI221XL U591 (.Y(n1266), 
	.C0(n682), 
	.B1(n465), 
	.B0(n1344), 
	.A1(n236), 
	.A0(n681));
   XNOR2X1 U592 (.Y(n681), 
	.B(block[66]), 
	.A(round_key[66]));
   AOI222X1 U593 (.Y(n682), 
	.C1(n684), 
	.C0(FE_OFN98_n232), 
	.B1(n683), 
	.B0(n96), 
	.A1(new_sboxw[2]), 
	.A0(n4));
   XNOR2X1 U594 (.Y(n683), 
	.B(n1395), 
	.A(round_key[66]));
   OAI221XL U595 (.Y(n1293), 
	.C0(n886), 
	.B1(n706), 
	.B0(n1341), 
	.A1(n108), 
	.A0(n885));
   XNOR2X1 U596 (.Y(n885), 
	.B(block[39]), 
	.A(round_key[39]));
   AOI222X1 U597 (.Y(n886), 
	.C1(n888), 
	.C0(FE_OFN97_n232), 
	.B1(n887), 
	.B0(n97), 
	.A1(new_sboxw[7]), 
	.A0(n16));
   XNOR2X1 U598 (.Y(n887), 
	.B(n1412), 
	.A(round_key[39]));
   OAI221XL U599 (.Y(n1327), 
	.C0(n1139), 
	.B1(n945), 
	.B0(n192), 
	.A1(n108), 
	.A0(FE_PHN5244_n1138));
   XNOR2X1 U600 (.Y(n1138), 
	.B(block[5]), 
	.A(round_key[5]));
   AOI222X1 U601 (.Y(n1139), 
	.C1(n1141), 
	.C0(FE_OFN97_n232), 
	.B1(n1140), 
	.B0(n96), 
	.A1(new_sboxw[5]), 
	.A0(n7));
   XNOR2X1 U602 (.Y(n1140), 
	.B(n191), 
	.A(round_key[5]));
   OAI221XL U603 (.Y(n1295), 
	.C0(n900), 
	.B1(n706), 
	.B0(n191), 
	.A1(n108), 
	.A0(n899));
   XNOR2X1 U604 (.Y(n899), 
	.B(block[37]), 
	.A(round_key[37]));
   AOI222X1 U605 (.Y(n900), 
	.C1(n902), 
	.C0(FE_OFN97_n232), 
	.B1(n901), 
	.B0(n97), 
	.A1(new_sboxw[5]), 
	.A0(n16));
   XNOR2X1 U606 (.Y(n901), 
	.B(n1352), 
	.A(round_key[37]));
   OAI221XL U607 (.Y(n1290), 
	.C0(n867), 
	.B1(n706), 
	.B0(n186), 
	.A1(n108), 
	.A0(FE_PHN5207_n866));
   XNOR2X1 U608 (.Y(n866), 
	.B(block[42]), 
	.A(round_key[42]));
   AOI222X1 U609 (.Y(n867), 
	.C1(n869), 
	.C0(FE_OFN98_n232), 
	.B1(n868), 
	.B0(n97), 
	.A1(new_sboxw[10]), 
	.A0(n16));
   XNOR2X1 U610 (.Y(n868), 
	.B(n1361), 
	.A(round_key[42]));
   OAI221XL U611 (.Y(n1219), 
	.C0(n340), 
	.B1(n230), 
	.B0(n1443), 
	.A1(n105), 
	.A0(n339));
   XNOR2X1 U612 (.Y(n339), 
	.B(block[114]), 
	.A(round_key[114]));
   AOI222X1 U613 (.Y(n340), 
	.C1(n342), 
	.C0(n232), 
	.B1(n341), 
	.B0(n96), 
	.A1(n13), 
	.A0(new_sboxw[18]));
   XNOR2X1 U614 (.Y(n341), 
	.B(n1441), 
	.A(round_key[114]));
   OAI221XL U615 (.Y(n1214), 
	.C0(n302), 
	.B1(n230), 
	.B0(n1415), 
	.A1(n107), 
	.A0(n301));
   XNOR2X1 U616 (.Y(n301), 
	.B(block[119]), 
	.A(round_key[119]));
   AOI222X1 U617 (.Y(n302), 
	.C1(n304), 
	.C0(FE_OFN97_n232), 
	.B1(n303), 
	.B0(n96), 
	.A1(n13), 
	.A0(new_sboxw[23]));
   XNOR2X1 U618 (.Y(n303), 
	.B(n1414), 
	.A(round_key[119]));
   OAI221XL U619 (.Y(n1235), 
	.C0(n450), 
	.B1(n230), 
	.B0(n1395), 
	.A1(n99), 
	.A0(n449));
   XNOR2X1 U620 (.Y(n449), 
	.B(block[98]), 
	.A(round_key[98]));
   AOI222X1 U621 (.Y(n450), 
	.C1(n452), 
	.C0(n232), 
	.B1(n451), 
	.B0(n96), 
	.A1(n12), 
	.A0(new_sboxw[2]));
   XNOR2X1 U622 (.Y(n451), 
	.B(n1454), 
	.A(round_key[98]));
   OAI221XL U623 (.Y(n1227), 
	.C0(n394), 
	.B1(n230), 
	.B0(n1361), 
	.A1(n99), 
	.A0(n393));
   XNOR2X1 U624 (.Y(n393), 
	.B(block[106]), 
	.A(round_key[106]));
   AOI222X1 U625 (.Y(n394), 
	.C1(n396), 
	.C0(n232), 
	.B1(n395), 
	.B0(n96), 
	.A1(n12), 
	.A0(new_sboxw[10]));
   XNOR2X1 U626 (.Y(n395), 
	.B(n186), 
	.A(round_key[106]));
   OAI221XL U627 (.Y(n1230), 
	.C0(n413), 
	.B1(n230), 
	.B0(n1357), 
	.A1(n99), 
	.A0(n412));
   XNOR2X1 U628 (.Y(n412), 
	.B(block[103]), 
	.A(round_key[103]));
   AOI222X1 U629 (.Y(n413), 
	.C1(n415), 
	.C0(FE_OFN97_n232), 
	.B1(n414), 
	.B0(n96), 
	.A1(n12), 
	.A0(new_sboxw[7]));
   XNOR2X1 U630 (.Y(n414), 
	.B(n1381), 
	.A(round_key[103]));
   OAI221XL U631 (.Y(n1222), 
	.C0(n361), 
	.B1(n230), 
	.B0(n1199), 
	.A1(n99), 
	.A0(n360));
   XNOR2X1 U632 (.Y(n360), 
	.B(block[111]), 
	.A(round_key[111]));
   AOI222X1 U633 (.Y(n361), 
	.C1(n363), 
	.C0(FE_OFN97_n232), 
	.B1(n362), 
	.B0(n38), 
	.A1(n13), 
	.A0(new_sboxw[15]));
   XNOR2X1 U634 (.Y(n362), 
	.B(n1356), 
	.A(round_key[111]));
   OAI221XL U635 (.Y(n1246), 
	.C0(n542), 
	.B1(n465), 
	.B0(n1411), 
	.A1(n106), 
	.A0(FE_PHN5134_n541));
   XNOR2X1 U636 (.Y(n541), 
	.B(block[86]), 
	.A(round_key[86]));
   AOI222X1 U637 (.Y(n542), 
	.C1(n544), 
	.C0(FE_OFN97_n232), 
	.B1(n543), 
	.B0(n96), 
	.A1(new_sboxw[22]), 
	.A0(n11));
   XNOR2X1 U638 (.Y(n543), 
	.B(n1409), 
	.A(round_key[86]));
   OAI221XL U639 (.Y(n1278), 
	.C0(n783), 
	.B1(n706), 
	.B0(n1409), 
	.A1(n236), 
	.A0(FE_PHN5150_n782));
   XNOR2X1 U640 (.Y(n782), 
	.B(block[54]), 
	.A(round_key[54]));
   AOI222X1 U641 (.Y(n783), 
	.C1(n785), 
	.C0(FE_OFN97_n232), 
	.B1(n784), 
	.B0(n97), 
	.A1(new_sboxw[22]), 
	.A0(n17));
   XNOR2X1 U642 (.Y(n784), 
	.B(n1408), 
	.A(round_key[54]));
   OAI221XL U643 (.Y(n1310), 
	.C0(n1022), 
	.B1(n945), 
	.B0(n1408), 
	.A1(n107), 
	.A0(FE_PHN5126_n1021));
   XNOR2X1 U644 (.Y(n1021), 
	.B(block[22]), 
	.A(round_key[22]));
   AOI222X1 U645 (.Y(n1022), 
	.C1(n1024), 
	.C0(FE_OFN97_n232), 
	.B1(n1023), 
	.B0(n83), 
	.A1(new_sboxw[22]), 
	.A0(n8));
   XNOR2X1 U646 (.Y(n1023), 
	.B(n1407), 
	.A(round_key[22]));
   OAI221XL U647 (.Y(n1318), 
	.C0(n1079), 
	.B1(n945), 
	.B0(n1378), 
	.A1(n107), 
	.A0(FE_PHN5144_n1078));
   XNOR2X1 U648 (.Y(n1078), 
	.B(block[14]), 
	.A(round_key[14]));
   AOI222X1 U649 (.Y(n1079), 
	.C1(n1081), 
	.C0(FE_OFN97_n232), 
	.B1(n1080), 
	.B0(n97), 
	.A1(new_sboxw[14]), 
	.A0(n8));
   XNOR2X1 U650 (.Y(n1080), 
	.B(n1367), 
	.A(round_key[14]));
   OAI221XL U651 (.Y(n1254), 
	.C0(n599), 
	.B1(n465), 
	.B0(n1367), 
	.A1(n106), 
	.A0(n598));
   XNOR2X1 U652 (.Y(n598), 
	.B(block[78]), 
	.A(round_key[78]));
   AOI222X1 U653 (.Y(n599), 
	.C1(n601), 
	.C0(FE_OFN97_n232), 
	.B1(n600), 
	.B0(n49), 
	.A1(new_sboxw[14]), 
	.A0(n11));
   XNOR2X1 U654 (.Y(n600), 
	.B(n1378), 
	.A(round_key[78]));
   OAI221XL U655 (.Y(n1262), 
	.C0(n652), 
	.B1(n465), 
	.B0(n1355), 
	.A1(n236), 
	.A0(FE_PHN5119_n651));
   XNOR2X1 U656 (.Y(n651), 
	.B(block[70]), 
	.A(round_key[70]));
   AOI222X1 U657 (.Y(n652), 
	.C1(n654), 
	.C0(FE_OFN97_n232), 
	.B1(n653), 
	.B0(n96), 
	.A1(new_sboxw[6]), 
	.A0(n4));
   XNOR2X1 U658 (.Y(n653), 
	.B(n1354), 
	.A(round_key[70]));
   OAI221XL U659 (.Y(n1286), 
	.C0(n840), 
	.B1(n706), 
	.B0(n1353), 
	.A1(n107), 
	.A0(n839));
   XNOR2X1 U660 (.Y(n839), 
	.B(block[46]), 
	.A(round_key[46]));
   AOI222X1 U661 (.Y(n840), 
	.C1(n842), 
	.C0(FE_OFN97_n232), 
	.B1(n841), 
	.B0(n97), 
	.A1(new_sboxw[14]), 
	.A0(n17));
   XNOR2X1 U662 (.Y(n841), 
	.B(n229), 
	.A(round_key[46]));
   OAI221XL U663 (.Y(n1326), 
	.C0(n1132), 
	.B1(n945), 
	.B0(n944), 
	.A1(n108), 
	.A0(FE_PHN5102_n1131));
   XNOR2X1 U664 (.Y(n1131), 
	.B(block[6]), 
	.A(round_key[6]));
   AOI222X1 U665 (.Y(n1132), 
	.C1(n1134), 
	.C0(FE_OFN97_n232), 
	.B1(n1133), 
	.B0(n96), 
	.A1(new_sboxw[6]), 
	.A0(n7));
   XNOR2X1 U666 (.Y(n1133), 
	.B(n705), 
	.A(round_key[6]));
   OAI221XL U667 (.Y(n1294), 
	.C0(n893), 
	.B1(n706), 
	.B0(n705), 
	.A1(n106), 
	.A0(FE_PHN5256_n892));
   XNOR2X1 U668 (.Y(n892), 
	.B(block[38]), 
	.A(round_key[38]));
   AOI222X1 U669 (.Y(n893), 
	.C1(n895), 
	.C0(FE_OFN97_n232), 
	.B1(n894), 
	.B0(n97), 
	.A1(new_sboxw[6]), 
	.A0(n16));
   XNOR2X1 U670 (.Y(n894), 
	.B(n1355), 
	.A(round_key[38]));
   OAI221XL U671 (.Y(n1324), 
	.C0(n1119), 
	.B1(n945), 
	.B0(n1425), 
	.A1(n108), 
	.A0(n1118));
   XNOR2X1 U672 (.Y(n1118), 
	.B(block[8]), 
	.A(round_key[8]));
   AOI222X1 U673 (.Y(n1119), 
	.C1(n1121), 
	.C0(FE_OFN98_n232), 
	.B1(n1120), 
	.B0(n96), 
	.A1(new_sboxw[8]), 
	.A0(n7));
   XNOR2X1 U674 (.Y(n1120), 
	.B(n1369), 
	.A(round_key[8]));
   OAI221XL U675 (.Y(n1236), 
	.C0(n457), 
	.B1(n230), 
	.B0(n1343), 
	.A1(n107), 
	.A0(n456));
   XNOR2X1 U676 (.Y(n456), 
	.B(block[97]), 
	.A(round_key[97]));
   AOI222X1 U677 (.Y(n457), 
	.C1(n459), 
	.C0(FE_OFN98_n232), 
	.B1(n458), 
	.B0(n96), 
	.A1(n12), 
	.A0(new_sboxw[1]));
   XNOR2X1 U678 (.Y(n458), 
	.B(n1394), 
	.A(round_key[97]));
   OAI221XL U679 (.Y(n1331), 
	.C0(n1169), 
	.B1(n945), 
	.B0(n1394), 
	.A1(n108), 
	.A0(n1168));
   XNOR2X1 U680 (.Y(n1168), 
	.B(block[1]), 
	.A(round_key[1]));
   AOI222X1 U681 (.Y(n1169), 
	.C1(n1171), 
	.C0(FE_OFN98_n232), 
	.B1(n1170), 
	.B0(n96), 
	.A1(new_sboxw[1]), 
	.A0(n7));
   XNOR2X1 U682 (.Y(n1170), 
	.B(n1453), 
	.A(round_key[1]));
   OAI221XL U683 (.Y(n1233), 
	.C0(n434), 
	.B1(n230), 
	.B0(n1364), 
	.A1(n106), 
	.A0(n433));
   XNOR2X1 U684 (.Y(n433), 
	.B(block[100]), 
	.A(round_key[100]));
   AOI222X1 U685 (.Y(n434), 
	.C1(n436), 
	.C0(FE_OFN98_n232), 
	.B1(n435), 
	.B0(n96), 
	.A1(n12), 
	.A0(new_sboxw[4]));
   XNOR2X1 U686 (.Y(n435), 
	.B(n189), 
	.A(round_key[100]));
   OAI221XL U687 (.Y(n1231), 
	.C0(n420), 
	.B1(n230), 
	.B0(n1354), 
	.A1(n99), 
	.A0(FE_PHN5075_n419));
   XNOR2X1 U688 (.Y(n419), 
	.B(block[102]), 
	.A(round_key[102]));
   AOI222X1 U689 (.Y(n420), 
	.C1(n422), 
	.C0(FE_OFN97_n232), 
	.B1(n421), 
	.B0(n96), 
	.A1(n12), 
	.A0(new_sboxw[6]));
   XNOR2X1 U690 (.Y(n421), 
	.B(n944), 
	.A(round_key[102]));
   OAI221XL U691 (.Y(n1232), 
	.C0(n427), 
	.B1(n230), 
	.B0(n1351), 
	.A1(n106), 
	.A0(FE_PHN5161_n426));
   XNOR2X1 U692 (.Y(n426), 
	.B(block[101]), 
	.A(round_key[101]));
   AOI222X1 U693 (.Y(n427), 
	.C1(n429), 
	.C0(FE_OFN97_n232), 
	.B1(n428), 
	.B0(n96), 
	.A1(n12), 
	.A0(new_sboxw[5]));
   XNOR2X1 U694 (.Y(n428), 
	.B(n192), 
	.A(round_key[101]));
   OAI221XL U695 (.Y(n1223), 
	.C0(n367), 
	.B1(n230), 
	.B0(n229), 
	.A1(n105), 
	.A0(FE_PHN5125_n366));
   XNOR2X1 U696 (.Y(n366), 
	.B(block[110]), 
	.A(round_key[110]));
   AOI222X1 U697 (.Y(n367), 
	.C1(n369), 
	.C0(FE_OFN97_n232), 
	.B1(n368), 
	.B0(n39), 
	.A1(n13), 
	.A0(new_sboxw[14]));
   XNOR2X1 U698 (.Y(n368), 
	.B(n1353), 
	.A(round_key[110]));
   OAI221XL U699 (.Y(n1224), 
	.C0(n373), 
	.B1(n230), 
	.B0(n190), 
	.A1(n107), 
	.A0(FE_PHN5148_n372));
   XNOR2X1 U700 (.Y(n372), 
	.B(block[109]), 
	.A(round_key[109]));
   AOI222X1 U701 (.Y(n373), 
	.C1(n375), 
	.C0(FE_OFN97_n232), 
	.B1(n374), 
	.B0(n39), 
	.A1(n13), 
	.A0(new_sboxw[13]));
   XNOR2X1 U702 (.Y(n374), 
	.B(n1350), 
	.A(round_key[109]));
   OAI221XL U703 (.Y(n1206), 
	.C0(n231), 
	.B1(n230), 
	.B0(n1417), 
	.A1(n139), 
	.A0(n1));
   AOI222X1 U704 (.Y(n231), 
	.C1(n235), 
	.C0(round_key[127]), 
	.B1(n169), 
	.B0(n234), 
	.A1(n233), 
	.A0(FE_OFN97_n232));
   OAI2BB2X1 U705 (.Y(n234), 
	.B1(FE_PHN157_n237), 
	.B0(n1417), 
	.A1N(block[127]), 
	.A0N(n110));
   OAI22X1 U706 (.Y(n235), 
	.B1(n30), 
	.B0(new_block[127]), 
	.A1(n105), 
	.A0(block[127]));
   OAI221XL U707 (.Y(n1207), 
	.C0(n242), 
	.B1(n230), 
	.B0(n1406), 
	.A1(n137), 
	.A0(n1));
   AOI222X1 U708 (.Y(n242), 
	.C1(n245), 
	.C0(round_key[126]), 
	.B1(n161), 
	.B0(n244), 
	.A1(n243), 
	.A0(FE_OFN97_n232));
   OAI2BB2X1 U709 (.Y(n244), 
	.B1(FE_PHN157_n237), 
	.B0(n1406), 
	.A1N(block[126]), 
	.A0N(n111));
   OAI22X1 U710 (.Y(n245), 
	.B1(n30), 
	.B0(new_block[126]), 
	.A1(n105), 
	.A0(block[126]));
   OAI221XL U711 (.Y(n1208), 
	.C0(n250), 
	.B1(n230), 
	.B0(n1405), 
	.A1(n138), 
	.A0(n1));
   AOI222X1 U712 (.Y(n250), 
	.C1(n253), 
	.C0(round_key[125]), 
	.B1(n157), 
	.B0(n252), 
	.A1(n251), 
	.A0(FE_OFN97_n232));
   OAI2BB2X1 U713 (.Y(n252), 
	.B1(FE_PHN157_n237), 
	.B0(n1405), 
	.A1N(block[125]), 
	.A0N(n113));
   OAI22X1 U714 (.Y(n253), 
	.B1(FE_PHN157_n237), 
	.B0(new_block[125]), 
	.A1(n105), 
	.A0(block[125]));
   OAI221XL U715 (.Y(n1323), 
	.C0(n1112), 
	.B1(n945), 
	.B0(n1370), 
	.A1(n108), 
	.A0(n1111));
   XNOR2X1 U716 (.Y(n1111), 
	.B(block[9]), 
	.A(round_key[9]));
   AOI222X1 U717 (.Y(n1112), 
	.C1(n1114), 
	.C0(FE_OFN98_n232), 
	.B1(n1113), 
	.B0(n96), 
	.A1(new_sboxw[9]), 
	.A0(n7));
   XNOR2X1 U718 (.Y(n1113), 
	.B(n1434), 
	.A(round_key[9]));
   OAI221XL U719 (.Y(n1328), 
	.C0(n1146), 
	.B1(n945), 
	.B0(n189), 
	.A1(n108), 
	.A0(n1145));
   XNOR2X1 U720 (.Y(n1145), 
	.B(block[4]), 
	.A(round_key[4]));
   AOI222X1 U721 (.Y(n1146), 
	.C1(n1148), 
	.C0(FE_OFN97_n232), 
	.B1(n1147), 
	.B0(n96), 
	.A1(new_sboxw[4]), 
	.A0(n7));
   XNOR2X1 U722 (.Y(n1147), 
	.B(n1347), 
	.A(round_key[4]));
   OAI221XL U723 (.Y(n1234), 
	.C0(n442), 
	.B1(n230), 
	.B0(n1382), 
	.A1(n106), 
	.A0(FE_PHN5110_n441));
   XNOR2X1 U724 (.Y(n441), 
	.B(block[99]), 
	.A(round_key[99]));
   AOI222X1 U725 (.Y(n442), 
	.C1(n444), 
	.C0(FE_OFN98_n232), 
	.B1(n443), 
	.B0(n96), 
	.A1(n12), 
	.A0(new_sboxw[3]));
   XNOR2X1 U726 (.Y(n443), 
	.B(n1452), 
	.A(round_key[99]));
   OAI221XL U727 (.Y(n1299), 
	.C0(n930), 
	.B1(n706), 
	.B0(n1453), 
	.A1(n107), 
	.A0(FE_PHN5233_n929));
   XNOR2X1 U728 (.Y(n929), 
	.B(block[33]), 
	.A(round_key[33]));
   AOI222X1 U729 (.Y(n930), 
	.C1(n932), 
	.C0(FE_OFN98_n232), 
	.B1(n931), 
	.B0(n97), 
	.A1(new_sboxw[1]), 
	.A0(n16));
   XNOR2X1 U730 (.Y(n931), 
	.B(n185), 
	.A(round_key[33]));
   OAI221XL U731 (.Y(n1288), 
	.C0(n852), 
	.B1(n706), 
	.B0(n1374), 
	.A1(n106), 
	.A0(n851));
   XNOR2X1 U732 (.Y(n851), 
	.B(block[44]), 
	.A(round_key[44]));
   AOI222X1 U733 (.Y(n852), 
	.C1(n854), 
	.C0(FE_OFN98_n232), 
	.B1(n853), 
	.B0(n97), 
	.A1(new_sboxw[12]), 
	.A0(n17));
   XNOR2X1 U734 (.Y(n853), 
	.B(n1346), 
	.A(round_key[44]));
   OAI221XL U735 (.Y(n1296), 
	.C0(n907), 
	.B1(n706), 
	.B0(n1347), 
	.A1(n106), 
	.A0(n906));
   XNOR2X1 U736 (.Y(n906), 
	.B(block[36]), 
	.A(round_key[36]));
   AOI222X1 U737 (.Y(n907), 
	.C1(n909), 
	.C0(FE_OFN98_n232), 
	.B1(n908), 
	.B0(n97), 
	.A1(new_sboxw[4]), 
	.A0(n16));
   XNOR2X1 U738 (.Y(n908), 
	.B(n1349), 
	.A(round_key[36]));
   OAI221XL U739 (.Y(n1329), 
	.C0(n1154), 
	.B1(n945), 
	.B0(n1452), 
	.A1(n108), 
	.A0(n1153));
   XNOR2X1 U740 (.Y(n1153), 
	.B(block[3]), 
	.A(round_key[3]));
   AOI222X1 U741 (.Y(n1154), 
	.C1(n1156), 
	.C0(FE_OFN98_n232), 
	.B1(n1155), 
	.B0(n96), 
	.A1(new_sboxw[3]), 
	.A0(n7));
   XNOR2X1 U742 (.Y(n1155), 
	.B(n188), 
	.A(round_key[3]));
   OAI221XL U743 (.Y(n1332), 
	.C0(n1177), 
	.B1(n945), 
	.B0(n1342), 
	.A1(n99), 
	.A0(n1176));
   XNOR2X1 U744 (.Y(n1176), 
	.B(block[0]), 
	.A(round_key[0]));
   AOI222X1 U745 (.Y(n1177), 
	.C1(n1179), 
	.C0(FE_OFN98_n232), 
	.B1(n1178), 
	.B0(n96), 
	.A1(new_sboxw[0]), 
	.A0(n7));
   OAI221XL U746 (.Y(n1229), 
	.C0(n407), 
	.B1(n230), 
	.B0(n1419), 
	.A1(n107), 
	.A0(n406));
   XNOR2X1 U747 (.Y(n406), 
	.B(block[104]), 
	.A(round_key[104]));
   AOI222X1 U748 (.Y(n407), 
	.C1(n409), 
	.C0(FE_OFN98_n232), 
	.B1(n408), 
	.B0(n96), 
	.A1(n12), 
	.A0(new_sboxw[8]));
   XNOR2X1 U749 (.Y(n408), 
	.B(n1420), 
	.A(round_key[104]));
   OAI221XL U750 (.Y(n1213), 
	.C0(n294), 
	.B1(n230), 
	.B0(n1418), 
	.A1(n143), 
	.A0(n1));
   AOI222X1 U751 (.Y(n294), 
	.C1(n297), 
	.C0(round_key[120]), 
	.B1(n165), 
	.B0(n296), 
	.A1(n295), 
	.A0(n232));
   OAI2BB2X1 U752 (.Y(n296), 
	.B1(FE_PHN157_n237), 
	.B0(n1418), 
	.A1N(block[120]), 
	.A0N(n113));
   OAI22X1 U753 (.Y(n297), 
	.B1(n30), 
	.B0(new_block[120]), 
	.A1(n105), 
	.A0(block[120]));
   OAI221XL U754 (.Y(n1239), 
	.C0(n482), 
	.B1(n465), 
	.B0(n1400), 
	.A1(n464), 
	.A0(n138));
   AOI222X1 U755 (.Y(n482), 
	.C1(n485), 
	.C0(round_key[93]), 
	.B1(n158), 
	.B0(n484), 
	.A1(n483), 
	.A0(FE_OFN97_n232));
   OAI2BB2X1 U756 (.Y(n484), 
	.B1(FE_PHN157_n237), 
	.B0(n1400), 
	.A1N(block[93]), 
	.A0N(n110));
   OAI22X1 U757 (.Y(n485), 
	.B1(n30), 
	.B0(new_block[93]), 
	.A1(n105), 
	.A0(block[93]));
   OAI221XL U758 (.Y(n1240), 
	.C0(n490), 
	.B1(n465), 
	.B0(n1399), 
	.A1(n464), 
	.A0(n140));
   AOI222X1 U759 (.Y(n490), 
	.C1(n493), 
	.C0(round_key[92]), 
	.B1(n154), 
	.B0(n492), 
	.A1(n491), 
	.A0(FE_OFN97_n232));
   OAI2BB2X1 U760 (.Y(n492), 
	.B1(FE_PHN157_n237), 
	.B0(n1399), 
	.A1N(block[92]), 
	.A0N(n114));
   OAI22X1 U761 (.Y(n493), 
	.B1(n30), 
	.B0(new_block[92]), 
	.A1(n105), 
	.A0(block[92]));
   OAI221XL U762 (.Y(n1285), 
	.C0(n834), 
	.B1(n706), 
	.B0(n1356), 
	.A1(n99), 
	.A0(n833));
   XNOR2X1 U763 (.Y(n833), 
	.B(block[47]), 
	.A(round_key[47]));
   AOI222X1 U764 (.Y(n834), 
	.C1(n836), 
	.C0(FE_OFN97_n232), 
	.B1(n835), 
	.B0(n97), 
	.A1(new_sboxw[15]), 
	.A0(n17));
   XNOR2X1 U765 (.Y(n835), 
	.B(n1199), 
	.A(round_key[47]));
   OAI221XL U766 (.Y(n1287), 
	.C0(n846), 
	.B1(n706), 
	.B0(n1350), 
	.A1(n107), 
	.A0(n845));
   XNOR2X1 U767 (.Y(n845), 
	.B(block[45]), 
	.A(round_key[45]));
   AOI222X1 U768 (.Y(n846), 
	.C1(n848), 
	.C0(FE_OFN97_n232), 
	.B1(n847), 
	.B0(n97), 
	.A1(new_sboxw[13]), 
	.A0(n17));
   XNOR2X1 U769 (.Y(n847), 
	.B(n190), 
	.A(round_key[45]));
   OAI221XL U770 (.Y(n1259), 
	.C0(n632), 
	.B1(n465), 
	.B0(n1434), 
	.A1(n236), 
	.A0(n631));
   XNOR2X1 U771 (.Y(n631), 
	.B(block[73]), 
	.A(round_key[73]));
   AOI222X1 U772 (.Y(n632), 
	.C1(n634), 
	.C0(FE_OFN98_n232), 
	.B1(n633), 
	.B0(n96), 
	.A1(new_sboxw[9]), 
	.A0(n4));
   XNOR2X1 U773 (.Y(n633), 
	.B(n1370), 
	.A(round_key[73]));
   OAI221XL U774 (.Y(n1255), 
	.C0(n605), 
	.B1(n465), 
	.B0(n1401), 
	.A1(n106), 
	.A0(n604));
   XNOR2X1 U775 (.Y(n604), 
	.B(block[77]), 
	.A(round_key[77]));
   AOI222X1 U776 (.Y(n605), 
	.C1(n607), 
	.C0(FE_OFN97_n232), 
	.B1(n606), 
	.B0(n50), 
	.A1(new_sboxw[13]), 
	.A0(n11));
   XNOR2X1 U777 (.Y(n606), 
	.B(n1366), 
	.A(round_key[77]));
   OAI221XL U778 (.Y(n1257), 
	.C0(n619), 
	.B1(n465), 
	.B0(n1396), 
	.A1(n106), 
	.A0(n618));
   XNOR2X1 U779 (.Y(n618), 
	.B(block[75]), 
	.A(round_key[75]));
   AOI222X1 U780 (.Y(n619), 
	.C1(n621), 
	.C0(FE_OFN98_n232), 
	.B1(n620), 
	.B0(n51), 
	.A1(new_sboxw[11]), 
	.A0(n4));
   XNOR2X1 U781 (.Y(n620), 
	.B(n1372), 
	.A(round_key[75]));
   OAI221XL U782 (.Y(n1265), 
	.C0(n674), 
	.B1(n465), 
	.B0(n1373), 
	.A1(n236), 
	.A0(n673));
   XNOR2X1 U783 (.Y(n673), 
	.B(block[67]), 
	.A(round_key[67]));
   AOI222X1 U784 (.Y(n674), 
	.C1(n676), 
	.C0(FE_OFN98_n232), 
	.B1(n675), 
	.B0(n96), 
	.A1(new_sboxw[3]), 
	.A0(n4));
   XNOR2X1 U785 (.Y(n675), 
	.B(n1382), 
	.A(round_key[67]));
   OAI221XL U786 (.Y(n1260), 
	.C0(n639), 
	.B1(n465), 
	.B0(n1369), 
	.A1(n236), 
	.A0(n638));
   XNOR2X1 U787 (.Y(n638), 
	.B(block[72]), 
	.A(round_key[72]));
   AOI222X1 U788 (.Y(n639), 
	.C1(n641), 
	.C0(FE_OFN98_n232), 
	.B1(n640), 
	.B0(n96), 
	.A1(new_sboxw[8]), 
	.A0(n4));
   XNOR2X1 U789 (.Y(n640), 
	.B(n1425), 
	.A(round_key[72]));
   OAI221XL U790 (.Y(n1256), 
	.C0(n611), 
	.B1(n465), 
	.B0(n1365), 
	.A1(n106), 
	.A0(n610));
   XNOR2X1 U791 (.Y(n610), 
	.B(block[76]), 
	.A(round_key[76]));
   AOI222X1 U792 (.Y(n611), 
	.C1(n613), 
	.C0(FE_OFN97_n232), 
	.B1(n612), 
	.B0(n50), 
	.A1(new_sboxw[12]), 
	.A0(n4));
   XNOR2X1 U793 (.Y(n612), 
	.B(n1348), 
	.A(round_key[76]));
   OAI221XL U794 (.Y(n1268), 
	.C0(n697), 
	.B1(n465), 
	.B0(n1359), 
	.A1(n236), 
	.A0(FE_PHN5109_n696));
   XNOR2X1 U795 (.Y(n696), 
	.B(block[64]), 
	.A(round_key[64]));
   AOI222X1 U796 (.Y(n697), 
	.C1(n699), 
	.C0(FE_OFN98_n232), 
	.B1(n698), 
	.B0(n96), 
	.A1(n4), 
	.A0(new_sboxw[0]));
   XNOR2X1 U797 (.Y(n698), 
	.B(n184), 
	.A(round_key[64]));
   OAI221XL U798 (.Y(n1264), 
	.C0(n666), 
	.B1(n465), 
	.B0(n1349), 
	.A1(n236), 
	.A0(n665));
   XNOR2X1 U799 (.Y(n665), 
	.B(block[68]), 
	.A(round_key[68]));
   AOI222X1 U800 (.Y(n666), 
	.C1(n668), 
	.C0(FE_OFN97_n232), 
	.B1(n667), 
	.B0(n96), 
	.A1(new_sboxw[4]), 
	.A0(n4));
   XNOR2X1 U801 (.Y(n667), 
	.B(n1364), 
	.A(round_key[68]));
   OAI221XL U802 (.Y(n1267), 
	.C0(n689), 
	.B1(n465), 
	.B0(n185), 
	.A1(n236), 
	.A0(n688));
   XNOR2X1 U803 (.Y(n688), 
	.B(block[65]), 
	.A(round_key[65]));
   AOI222X1 U804 (.Y(n689), 
	.C1(n691), 
	.C0(FE_OFN98_n232), 
	.B1(n690), 
	.B0(n96), 
	.A1(new_sboxw[1]), 
	.A0(n4));
   XNOR2X1 U805 (.Y(n690), 
	.B(n1343), 
	.A(round_key[65]));
   OAI221XL U806 (.Y(n1301), 
	.C0(n946), 
	.B1(n945), 
	.B0(n1380), 
	.A1(n3), 
	.A0(n139));
   AOI222X1 U807 (.Y(n946), 
	.C1(n949), 
	.C0(round_key[31]), 
	.B1(n172), 
	.B0(n948), 
	.A1(n947), 
	.A0(FE_OFN97_n232));
   OAI2BB2X1 U808 (.Y(n948), 
	.B1(FE_PHN157_n237), 
	.B0(n1380), 
	.A1N(block[31]), 
	.A0N(n114));
   OAI22X1 U809 (.Y(n949), 
	.B1(FE_PHN157_n237), 
	.B0(new_block[31]), 
	.A1(n105), 
	.A0(block[31]));
   OAI221XL U810 (.Y(n1302), 
	.C0(n954), 
	.B1(n945), 
	.B0(n1377), 
	.A1(n3), 
	.A0(n137));
   AOI222X1 U811 (.Y(n954), 
	.C1(n957), 
	.C0(round_key[30]), 
	.B1(n164), 
	.B0(n956), 
	.A1(n955), 
	.A0(FE_OFN97_n232));
   OAI2BB2X1 U812 (.Y(n956), 
	.B1(FE_PHN157_n237), 
	.B0(n1377), 
	.A1N(block[30]), 
	.A0N(n114));
   OAI22X1 U813 (.Y(n957), 
	.B1(FE_PHN157_n237), 
	.B0(new_block[30]), 
	.A1(n105), 
	.A0(block[30]));
   OAI221XL U814 (.Y(n1303), 
	.C0(n962), 
	.B1(n945), 
	.B0(n1376), 
	.A1(n3), 
	.A0(n138));
   AOI222X1 U815 (.Y(n962), 
	.C1(n965), 
	.C0(round_key[29]), 
	.B1(n160), 
	.B0(n964), 
	.A1(n963), 
	.A0(FE_OFN97_n232));
   OAI2BB2X1 U816 (.Y(n964), 
	.B1(FE_PHN157_n237), 
	.B0(n1376), 
	.A1N(block[29]), 
	.A0N(n114));
   OAI22X1 U817 (.Y(n965), 
	.B1(FE_PHN157_n237), 
	.B0(new_block[29]), 
	.A1(n105), 
	.A0(block[29]));
   OAI221XL U818 (.Y(n1315), 
	.C0(n1059), 
	.B1(n945), 
	.B0(n1436), 
	.A1(n107), 
	.A0(n1058));
   XNOR2X1 U819 (.Y(n1058), 
	.B(block[17]), 
	.A(round_key[17]));
   AOI222X1 U820 (.Y(n1059), 
	.C1(n1061), 
	.C0(n232), 
	.B1(n1060), 
	.B0(n83), 
	.A1(new_sboxw[17]), 
	.A0(n8));
   XNOR2X1 U821 (.Y(n1060), 
	.B(n1432), 
	.A(round_key[17]));
   OAI221XL U822 (.Y(n1311), 
	.C0(n1029), 
	.B1(n945), 
	.B0(n1402), 
	.A1(n107), 
	.A0(FE_PHN5167_n1028));
   XNOR2X1 U823 (.Y(n1028), 
	.B(block[21]), 
	.A(round_key[21]));
   AOI222X1 U824 (.Y(n1029), 
	.C1(n1031), 
	.C0(FE_OFN97_n232), 
	.B1(n1030), 
	.B0(n83), 
	.A1(new_sboxw[21]), 
	.A0(n8));
   XNOR2X1 U825 (.Y(n1030), 
	.B(n1375), 
	.A(round_key[21]));
   OAI221XL U826 (.Y(n1312), 
	.C0(n1036), 
	.B1(n945), 
	.B0(n1387), 
	.A1(n107), 
	.A0(FE_PHN5127_n1035));
   XNOR2X1 U827 (.Y(n1035), 
	.B(block[20]), 
	.A(round_key[20]));
   AOI222X1 U828 (.Y(n1036), 
	.C1(n1038), 
	.C0(FE_OFN97_n232), 
	.B1(n1037), 
	.B0(n83), 
	.A1(new_sboxw[20]), 
	.A0(n8));
   XNOR2X1 U829 (.Y(n1037), 
	.B(n1385), 
	.A(round_key[20]));
   OAI221XL U830 (.Y(n1317), 
	.C0(n1073), 
	.B1(n945), 
	.B0(n1368), 
	.A1(n107), 
	.A0(FE_PHN5168_n1072));
   XNOR2X1 U831 (.Y(n1072), 
	.B(block[15]), 
	.A(round_key[15]));
   AOI222X1 U832 (.Y(n1073), 
	.C1(n1075), 
	.C0(FE_OFN97_n232), 
	.B1(n1074), 
	.B0(n97), 
	.A1(new_sboxw[15]), 
	.A0(n8));
   XNOR2X1 U833 (.Y(n1074), 
	.B(n1379), 
	.A(round_key[15]));
   OAI221XL U834 (.Y(n1319), 
	.C0(n1085), 
	.B1(n945), 
	.B0(n1366), 
	.A1(n107), 
	.A0(n1084));
   XNOR2X1 U835 (.Y(n1084), 
	.B(block[13]), 
	.A(round_key[13]));
   AOI222X1 U836 (.Y(n1085), 
	.C1(n1087), 
	.C0(FE_OFN97_n232), 
	.B1(n1086), 
	.B0(n97), 
	.A1(new_sboxw[13]), 
	.A0(n8));
   XNOR2X1 U837 (.Y(n1086), 
	.B(n1401), 
	.A(round_key[13]));
   OAI221XL U838 (.Y(n1220), 
	.C0(n347), 
	.B1(n230), 
	.B0(n1432), 
	.A1(n106), 
	.A0(n346));
   XNOR2X1 U839 (.Y(n346), 
	.B(block[113]), 
	.A(round_key[113]));
   AOI222X1 U840 (.Y(n347), 
	.C1(n349), 
	.C0(n232), 
	.B1(n348), 
	.B0(n96), 
	.A1(n13), 
	.A0(new_sboxw[17]));
   XNOR2X1 U841 (.Y(n348), 
	.B(n1430), 
	.A(round_key[113]));
   OAI221XL U842 (.Y(n1215), 
	.C0(n310), 
	.B1(n230), 
	.B0(n1407), 
	.A1(n105), 
	.A0(FE_PHN5142_n309));
   XNOR2X1 U843 (.Y(n309), 
	.B(block[118]), 
	.A(round_key[118]));
   AOI222X1 U844 (.Y(n310), 
	.C1(n312), 
	.C0(FE_OFN97_n232), 
	.B1(n311), 
	.B0(n96), 
	.A1(n13), 
	.A0(new_sboxw[22]));
   XNOR2X1 U845 (.Y(n311), 
	.B(n1411), 
	.A(round_key[118]));
   OAI221XL U846 (.Y(n1217), 
	.C0(n324), 
	.B1(n230), 
	.B0(n1385), 
	.A1(n105), 
	.A0(FE_PHN5221_n323));
   XNOR2X1 U847 (.Y(n323), 
	.B(block[116]), 
	.A(round_key[116]));
   AOI222X1 U848 (.Y(n324), 
	.C1(n326), 
	.C0(FE_OFN97_n232), 
	.B1(n325), 
	.B0(n96), 
	.A1(n13), 
	.A0(new_sboxw[20]));
   XNOR2X1 U849 (.Y(n325), 
	.B(n1363), 
	.A(round_key[116]));
   OAI221XL U850 (.Y(n1216), 
	.C0(n317), 
	.B1(n230), 
	.B0(n1375), 
	.A1(n99), 
	.A0(FE_PHN5206_n316));
   XNOR2X1 U851 (.Y(n316), 
	.B(block[117]), 
	.A(round_key[117]));
   AOI222X1 U852 (.Y(n317), 
	.C1(n319), 
	.C0(FE_OFN97_n232), 
	.B1(n318), 
	.B0(n96), 
	.A1(n13), 
	.A0(new_sboxw[21]));
   XNOR2X1 U853 (.Y(n318), 
	.B(n1404), 
	.A(round_key[117]));
   OAI221XL U854 (.Y(n1211), 
	.C0(n277), 
	.B1(n230), 
	.B0(n1442), 
	.A1(n141), 
	.A0(n1));
   AOI222X1 U855 (.Y(n277), 
	.C1(n280), 
	.C0(round_key[122]), 
	.B1(n145), 
	.B0(n279), 
	.A1(n278), 
	.A0(n232));
   OAI2BB2X1 U856 (.Y(n279), 
	.B1(FE_PHN157_n237), 
	.B0(n1442), 
	.A1N(block[122]), 
	.A0N(n113));
   OAI22X1 U857 (.Y(n280), 
	.B1(FE_PHN157_n237), 
	.B0(new_block[122]), 
	.A1(n105), 
	.A0(block[122]));
   OAI221XL U858 (.Y(n1212), 
	.C0(n285), 
	.B1(n230), 
	.B0(n1431), 
	.A1(n142), 
	.A0(n1));
   AOI222X1 U859 (.Y(n285), 
	.C1(n288), 
	.C0(round_key[121]), 
	.B1(n133), 
	.B0(n287), 
	.A1(n286), 
	.A0(n232));
   OAI2BB2X1 U860 (.Y(n287), 
	.B1(FE_PHN157_n237), 
	.B0(n1431), 
	.A1N(block[121]), 
	.A0N(n113));
   OAI22X1 U861 (.Y(n288), 
	.B1(FE_PHN157_n237), 
	.B0(new_block[121]), 
	.A1(n105), 
	.A0(block[121]));
   OAI221XL U862 (.Y(n1209), 
	.C0(n258), 
	.B1(n230), 
	.B0(n1384), 
	.A1(n140), 
	.A0(n1));
   AOI222X1 U863 (.Y(n258), 
	.C1(n261), 
	.C0(round_key[124]), 
	.B1(n153), 
	.B0(n260), 
	.A1(n259), 
	.A0(FE_OFN97_n232));
   OAI2BB2X1 U864 (.Y(n260), 
	.B1(FE_PHN157_n237), 
	.B0(n1384), 
	.A1N(block[124]), 
	.A0N(n113));
   OAI22X1 U865 (.Y(n261), 
	.B1(FE_PHN157_n237), 
	.B0(new_block[124]), 
	.A1(n105), 
	.A0(block[124]));
   OAI221XL U866 (.Y(n1228), 
	.C0(n400), 
	.B1(n230), 
	.B0(n1433), 
	.A1(n106), 
	.A0(n399));
   XNOR2X1 U867 (.Y(n399), 
	.B(block[105]), 
	.A(round_key[105]));
   AOI222X1 U868 (.Y(n400), 
	.C1(n402), 
	.C0(FE_OFN98_n232), 
	.B1(n401), 
	.B0(n96), 
	.A1(n12), 
	.A0(new_sboxw[9]));
   XNOR2X1 U869 (.Y(n401), 
	.B(n1360), 
	.A(round_key[105]));
   OAI221XL U870 (.Y(n1225), 
	.C0(n379), 
	.B1(n230), 
	.B0(n1346), 
	.A1(n105), 
	.A0(FE_PHN5132_n378));
   XNOR2X1 U871 (.Y(n378), 
	.B(block[108]), 
	.A(round_key[108]));
   AOI222X1 U872 (.Y(n379), 
	.C1(n381), 
	.C0(FE_OFN97_n232), 
	.B1(n380), 
	.B0(n39), 
	.A1(n13), 
	.A0(new_sboxw[12]));
   XNOR2X1 U873 (.Y(n380), 
	.B(n1374), 
	.A(round_key[108]));
   OAI221XL U874 (.Y(n1238), 
	.C0(n474), 
	.B1(n465), 
	.B0(n1410), 
	.A1(n464), 
	.A0(n137));
   AOI222X1 U875 (.Y(n474), 
	.C1(n477), 
	.C0(round_key[94]), 
	.B1(n162), 
	.B0(n476), 
	.A1(n475), 
	.A0(FE_OFN97_n232));
   OAI2BB2X1 U876 (.Y(n476), 
	.B1(FE_PHN157_n237), 
	.B0(n1410), 
	.A1N(block[94]), 
	.A0N(n110));
   OAI22X1 U877 (.Y(n477), 
	.B1(n30), 
	.B0(new_block[94]), 
	.A1(n105), 
	.A0(block[94]));
   OAI221XL U878 (.Y(n1275), 
	.C0(n758), 
	.B1(n706), 
	.B0(n1437), 
	.A1(n2), 
	.A0(n142));
   AOI222X1 U879 (.Y(n758), 
	.C1(n761), 
	.C0(round_key[57]), 
	.B1(n135), 
	.B0(n760), 
	.A1(n759), 
	.A0(FE_OFN98_n232));
   OAI2BB2X1 U880 (.Y(n760), 
	.B1(FE_PHN157_n237), 
	.B0(n1437), 
	.A1N(block[57]), 
	.A0N(n114));
   OAI22X1 U881 (.Y(n761), 
	.B1(FE_PHN157_n237), 
	.B0(new_block[57]), 
	.A1(n105), 
	.A0(block[57]));
   OAI221XL U882 (.Y(n1270), 
	.C0(n715), 
	.B1(n706), 
	.B0(n1390), 
	.A1(n2), 
	.A0(n137));
   AOI222X1 U883 (.Y(n715), 
	.C1(n718), 
	.C0(round_key[62]), 
	.B1(n163), 
	.B0(n717), 
	.A1(n716), 
	.A0(FE_OFN97_n232));
   OAI2BB2X1 U884 (.Y(n717), 
	.B1(FE_PHN157_n237), 
	.B0(n1390), 
	.A1N(block[62]), 
	.A0N(n114));
   OAI22X1 U885 (.Y(n718), 
	.B1(n30), 
	.B0(new_block[62]), 
	.A1(n105), 
	.A0(block[62]));
   OAI221XL U886 (.Y(n1271), 
	.C0(n723), 
	.B1(n706), 
	.B0(n1389), 
	.A1(n2), 
	.A0(n138));
   AOI222X1 U887 (.Y(n723), 
	.C1(n726), 
	.C0(round_key[61]), 
	.B1(n159), 
	.B0(n725), 
	.A1(n724), 
	.A0(FE_OFN97_n232));
   OAI2BB2X1 U888 (.Y(n725), 
	.B1(FE_PHN157_n237), 
	.B0(n1389), 
	.A1N(block[61]), 
	.A0N(n114));
   OAI22X1 U889 (.Y(n726), 
	.B1(FE_PHN157_n237), 
	.B0(new_block[61]), 
	.A1(n105), 
	.A0(block[61]));
   OAI221XL U890 (.Y(n1272), 
	.C0(n731), 
	.B1(n706), 
	.B0(n1388), 
	.A1(n2), 
	.A0(n140));
   AOI222X1 U891 (.Y(n731), 
	.C1(n734), 
	.C0(round_key[60]), 
	.B1(n155), 
	.B0(n733), 
	.A1(n732), 
	.A0(FE_OFN97_n232));
   OAI2BB2X1 U892 (.Y(n733), 
	.B1(FE_PHN157_n237), 
	.B0(n1388), 
	.A1N(block[60]), 
	.A0N(n111));
   OAI22X1 U893 (.Y(n734), 
	.B1(FE_PHN157_n237), 
	.B0(new_block[60]), 
	.A1(n105), 
	.A0(block[60]));
   OAI221XL U894 (.Y(n1308), 
	.C0(n1006), 
	.B1(n945), 
	.B0(n1422), 
	.A1(n3), 
	.A0(n143));
   AOI222X1 U895 (.Y(n1006), 
	.C1(n1009), 
	.C0(round_key[24]), 
	.B1(n168), 
	.B0(n1008), 
	.A1(n1007), 
	.A0(n232));
   OAI2BB2X1 U896 (.Y(n1008), 
	.B1(FE_PHN157_n237), 
	.B0(n1422), 
	.A1N(block[24]), 
	.A0N(n111));
   OAI22X1 U897 (.Y(n1009), 
	.B1(FE_PHN157_n237), 
	.B0(new_block[24]), 
	.A1(n105), 
	.A0(block[24]));
   OAI221XL U898 (.Y(n1291), 
	.C0(n873), 
	.B1(n706), 
	.B0(n1360), 
	.A1(n106), 
	.A0(n872));
   XNOR2X1 U899 (.Y(n872), 
	.B(block[41]), 
	.A(round_key[41]));
   AOI222X1 U900 (.Y(n873), 
	.C1(n875), 
	.C0(FE_OFN98_n232), 
	.B1(n874), 
	.B0(n97), 
	.A1(new_sboxw[9]), 
	.A0(n16));
   XNOR2X1 U901 (.Y(n874), 
	.B(n1433), 
	.A(round_key[41]));
   OAI221XL U902 (.Y(n1300), 
	.C0(n938), 
	.B1(n706), 
	.B0(n1393), 
	.A1(n107), 
	.A0(n937));
   XNOR2X1 U903 (.Y(n937), 
	.B(block[32]), 
	.A(round_key[32]));
   AOI222X1 U904 (.Y(n938), 
	.C1(n940), 
	.C0(FE_OFN98_n232), 
	.B1(n939), 
	.B0(n97), 
	.A1(new_sboxw[0]), 
	.A0(n16));
   XNOR2X1 U905 (.Y(n939), 
	.B(n1359), 
	.A(round_key[32]));
   OAI221XL U906 (.Y(n1269), 
	.C0(n707), 
	.B1(n706), 
	.B0(n1391), 
	.A1(n2), 
	.A0(n139));
   AOI222X1 U907 (.Y(n707), 
	.C1(n710), 
	.C0(round_key[63]), 
	.B1(n171), 
	.B0(n709), 
	.A1(n708), 
	.A0(FE_OFN97_n232));
   OAI2BB2X1 U908 (.Y(n709), 
	.B1(FE_PHN157_n237), 
	.B0(n1391), 
	.A1N(block[63]), 
	.A0N(n114));
   OAI22X1 U909 (.Y(n710), 
	.B1(n30), 
	.B0(new_block[63]), 
	.A1(n105), 
	.A0(block[63]));
   OAI221XL U910 (.Y(n1297), 
	.C0(n915), 
	.B1(n706), 
	.B0(n188), 
	.A1(n107), 
	.A0(n914));
   XNOR2X1 U911 (.Y(n914), 
	.B(block[35]), 
	.A(round_key[35]));
   AOI222X1 U912 (.Y(n915), 
	.C1(n917), 
	.C0(FE_OFN98_n232), 
	.B1(n916), 
	.B0(n97), 
	.A1(new_sboxw[3]), 
	.A0(n16));
   XNOR2X1 U913 (.Y(n916), 
	.B(n1373), 
	.A(round_key[35]));
   OAI221XL U914 (.Y(n1333), 
	.C0(n1184), 
	.B1(n230), 
	.B0(n184), 
	.A1(n99), 
	.A0(n1183));
   XNOR2X1 U915 (.Y(n1183), 
	.B(block[96]), 
	.A(round_key[96]));
   AOI222X1 U916 (.Y(n1184), 
	.C1(n1186), 
	.C0(FE_OFN98_n232), 
	.B1(n1185), 
	.B0(n35), 
	.A1(n12), 
	.A0(new_sboxw[0]));
   XNOR2X1 U917 (.Y(n1185), 
	.B(n1342), 
	.A(round_key[96]));
   OAI221XL U918 (.Y(n1237), 
	.C0(n466), 
	.B1(n465), 
	.B0(n1358), 
	.A1(n464), 
	.A0(n139));
   AOI222X1 U919 (.Y(n466), 
	.C1(n469), 
	.C0(round_key[95]), 
	.B1(n170), 
	.B0(n468), 
	.A1(n467), 
	.A0(FE_OFN97_n232));
   OAI2BB2X1 U920 (.Y(n468), 
	.B1(FE_PHN157_n237), 
	.B0(n1358), 
	.A1N(block[95]), 
	.A0N(n114));
   OAI22X1 U921 (.Y(n469), 
	.B1(FE_PHN157_n237), 
	.B0(new_block[95]), 
	.A1(n105), 
	.A0(block[95]));
   OAI221XL U922 (.Y(n1306), 
	.C0(n989), 
	.B1(n945), 
	.B0(n1444), 
	.A1(n3), 
	.A0(n141));
   AOI222X1 U923 (.Y(n989), 
	.C1(n992), 
	.C0(round_key[26]), 
	.B1(n148), 
	.B0(n991), 
	.A1(n990), 
	.A0(n232));
   OAI2BB2X1 U924 (.Y(n991), 
	.B1(FE_PHN157_n237), 
	.B0(n1444), 
	.A1N(block[26]), 
	.A0N(n114));
   OAI22X1 U925 (.Y(n992), 
	.B1(FE_PHN157_n237), 
	.B0(new_block[26]), 
	.A1(n105), 
	.A0(block[26]));
   OAI221XL U926 (.Y(n1307), 
	.C0(n997), 
	.B1(n945), 
	.B0(n1435), 
	.A1(n3), 
	.A0(n142));
   AOI222X1 U927 (.Y(n997), 
	.C1(n1000), 
	.C0(round_key[25]), 
	.B1(n136), 
	.B0(n999), 
	.A1(n998), 
	.A0(n232));
   OAI2BB2X1 U928 (.Y(n999), 
	.B1(FE_PHN157_n237), 
	.B0(n1435), 
	.A1N(block[25]), 
	.A0N(n110));
   OAI22X1 U929 (.Y(n1000), 
	.B1(FE_PHN157_n237), 
	.B0(new_block[25]), 
	.A1(n105), 
	.A0(block[25]));
   OAI221XL U930 (.Y(n1304), 
	.C0(n970), 
	.B1(n945), 
	.B0(n1386), 
	.A1(n3), 
	.A0(n140));
   AOI222X1 U931 (.Y(n970), 
	.C1(n973), 
	.C0(round_key[28]), 
	.B1(n156), 
	.B0(n972), 
	.A1(n971), 
	.A0(FE_OFN97_n232));
   OAI2BB2X1 U932 (.Y(n972), 
	.B1(FE_PHN157_n237), 
	.B0(n1386), 
	.A1N(block[28]), 
	.A0N(n114));
   OAI22X1 U933 (.Y(n973), 
	.B1(FE_PHN157_n237), 
	.B0(new_block[28]), 
	.A1(n105), 
	.A0(block[28]));
   OAI221XL U934 (.Y(n1283), 
	.C0(n820), 
	.B1(n706), 
	.B0(n1428), 
	.A1(n106), 
	.A0(n819));
   XNOR2X1 U935 (.Y(n819), 
	.B(block[49]), 
	.A(round_key[49]));
   AOI222X1 U936 (.Y(n820), 
	.C1(n822), 
	.C0(FE_OFN98_n232), 
	.B1(n821), 
	.B0(n83), 
	.A1(new_sboxw[17]), 
	.A0(n17));
   XNOR2X1 U937 (.Y(n821), 
	.B(n1436), 
	.A(round_key[49]));
   OAI221XL U938 (.Y(n1279), 
	.C0(n790), 
	.B1(n706), 
	.B0(n1403), 
	.A1(n236), 
	.A0(n789));
   XNOR2X1 U939 (.Y(n789), 
	.B(block[53]), 
	.A(round_key[53]));
   AOI222X1 U940 (.Y(n790), 
	.C1(n792), 
	.C0(FE_OFN97_n232), 
	.B1(n791), 
	.B0(n97), 
	.A1(new_sboxw[21]), 
	.A0(n17));
   XNOR2X1 U941 (.Y(n791), 
	.B(n1402), 
	.A(round_key[53]));
   OAI221XL U942 (.Y(n1280), 
	.C0(n797), 
	.B1(n706), 
	.B0(n1398), 
	.A1(n236), 
	.A0(n796));
   XNOR2X1 U943 (.Y(n796), 
	.B(block[52]), 
	.A(round_key[52]));
   AOI222X1 U944 (.Y(n797), 
	.C1(n799), 
	.C0(FE_OFN97_n232), 
	.B1(n798), 
	.B0(n83), 
	.A1(new_sboxw[20]), 
	.A0(n17));
   XNOR2X1 U945 (.Y(n798), 
	.B(n1387), 
	.A(round_key[52]));
   OAI221XL U946 (.Y(n1241), 
	.C0(n500), 
	.B1(n465), 
	.B0(n1449), 
	.A1(n464), 
	.A0(n144));
   AOI222X1 U947 (.Y(n500), 
	.C1(n503), 
	.C0(round_key[91]), 
	.B1(n150), 
	.B0(n502), 
	.A1(n501), 
	.A0(FE_OFN98_n232));
   OAI2BB2X1 U948 (.Y(n502), 
	.B1(FE_PHN157_n237), 
	.B0(n1449), 
	.A1N(block[91]), 
	.A0N(n113));
   OAI22X1 U949 (.Y(n503), 
	.B1(n30), 
	.B0(new_block[91]), 
	.A1(n105), 
	.A0(block[91]));
   OAI221XL U950 (.Y(n1244), 
	.C0(n526), 
	.B1(n465), 
	.B0(n1426), 
	.A1(n464), 
	.A0(n143));
   AOI222X1 U951 (.Y(n526), 
	.C1(n529), 
	.C0(round_key[88]), 
	.B1(n166), 
	.B0(n528), 
	.A1(n527), 
	.A0(FE_OFN98_n232));
   OAI2BB2X1 U952 (.Y(n528), 
	.B1(FE_PHN157_n237), 
	.B0(n1426), 
	.A1N(block[88]), 
	.A0N(n114));
   OAI22X1 U953 (.Y(n529), 
	.B1(n30), 
	.B0(new_block[88]), 
	.A1(n105), 
	.A0(block[88]));
   OAI221XL U954 (.Y(n1273), 
	.C0(n741), 
	.B1(n706), 
	.B0(n1450), 
	.A1(n2), 
	.A0(n144));
   AOI222X1 U955 (.Y(n741), 
	.C1(n744), 
	.C0(round_key[59]), 
	.B1(n151), 
	.B0(n743), 
	.A1(n742), 
	.A0(FE_OFN98_n232));
   OAI2BB2X1 U956 (.Y(n743), 
	.B1(FE_PHN157_n237), 
	.B0(n1450), 
	.A1N(block[59]), 
	.A0N(n110));
   OAI22X1 U957 (.Y(n744), 
	.B1(FE_PHN157_n237), 
	.B0(new_block[59]), 
	.A1(n105), 
	.A0(block[59]));
   OAI221XL U958 (.Y(n1274), 
	.C0(n750), 
	.B1(n706), 
	.B0(n1438), 
	.A1(n2), 
	.A0(n141));
   AOI222X1 U959 (.Y(n750), 
	.C1(n753), 
	.C0(round_key[58]), 
	.B1(n147), 
	.B0(n752), 
	.A1(n751), 
	.A0(FE_OFN98_n232));
   OAI2BB2X1 U960 (.Y(n752), 
	.B1(FE_PHN157_n237), 
	.B0(n1438), 
	.A1N(block[58]), 
	.A0N(n110));
   OAI22X1 U961 (.Y(n753), 
	.B1(FE_PHN157_n237), 
	.B0(new_block[58]), 
	.A1(n105), 
	.A0(block[58]));
   OAI221XL U962 (.Y(n1276), 
	.C0(n767), 
	.B1(n706), 
	.B0(n1392), 
	.A1(n2), 
	.A0(n143));
   AOI222X1 U963 (.Y(n767), 
	.C1(n770), 
	.C0(round_key[56]), 
	.B1(n167), 
	.B0(n769), 
	.A1(n768), 
	.A0(FE_OFN98_n232));
   OAI2BB2X1 U964 (.Y(n769), 
	.B1(FE_PHN157_n237), 
	.B0(n1392), 
	.A1N(block[56]), 
	.A0N(n114));
   OAI22X1 U965 (.Y(n770), 
	.B1(FE_PHN157_n237), 
	.B0(new_block[56]), 
	.A1(n105), 
	.A0(block[56]));
   OAI221XL U966 (.Y(n1210), 
	.C0(n268), 
	.B1(n230), 
	.B0(n1446), 
	.A1(n144), 
	.A0(n1));
   AOI222X1 U967 (.Y(n268), 
	.C1(n271), 
	.C0(round_key[123]), 
	.B1(n149), 
	.B0(n270), 
	.A1(n269), 
	.A0(FE_OFN97_n232));
   OAI2BB2X1 U968 (.Y(n270), 
	.B1(FE_PHN157_n237), 
	.B0(n1446), 
	.A1N(block[123]), 
	.A0N(n113));
   OAI22X1 U969 (.Y(n271), 
	.B1(n30), 
	.B0(new_block[123]), 
	.A1(n105), 
	.A0(block[123]));
   OAI221XL U970 (.Y(n1251), 
	.C0(n579), 
	.B1(n465), 
	.B0(n1430), 
	.A1(n106), 
	.A0(n578));
   XNOR2X1 U971 (.Y(n578), 
	.B(block[81]), 
	.A(round_key[81]));
   AOI222X1 U972 (.Y(n579), 
	.C1(n581), 
	.C0(FE_OFN98_n232), 
	.B1(n580), 
	.B0(n48), 
	.A1(new_sboxw[17]), 
	.A0(n11));
   XNOR2X1 U973 (.Y(n580), 
	.B(n1428), 
	.A(round_key[81]));
   OAI221XL U974 (.Y(n1252), 
	.C0(n587), 
	.B1(n465), 
	.B0(n1427), 
	.A1(n106), 
	.A0(n586));
   XNOR2X1 U975 (.Y(n586), 
	.B(block[80]), 
	.A(round_key[80]));
   AOI222X1 U976 (.Y(n587), 
	.C1(n589), 
	.C0(FE_OFN98_n232), 
	.B1(n588), 
	.B0(n48), 
	.A1(new_sboxw[16]), 
	.A0(n11));
   XNOR2X1 U977 (.Y(n588), 
	.B(n1424), 
	.A(round_key[80]));
   OAI221XL U978 (.Y(n1247), 
	.C0(n549), 
	.B1(n465), 
	.B0(n1404), 
	.A1(n106), 
	.A0(FE_PHN5146_n548));
   XNOR2X1 U979 (.Y(n548), 
	.B(block[85]), 
	.A(round_key[85]));
   AOI222X1 U980 (.Y(n549), 
	.C1(n551), 
	.C0(FE_OFN97_n232), 
	.B1(n550), 
	.B0(n46), 
	.A1(new_sboxw[21]), 
	.A0(n11));
   XNOR2X1 U981 (.Y(n550), 
	.B(n1403), 
	.A(round_key[85]));
   OAI221XL U982 (.Y(n1249), 
	.C0(n564), 
	.B1(n465), 
	.B0(n1383), 
	.A1(n106), 
	.A0(FE_PHN5165_n563));
   XNOR2X1 U983 (.Y(n563), 
	.B(block[83]), 
	.A(round_key[83]));
   AOI222X1 U984 (.Y(n564), 
	.C1(n566), 
	.C0(FE_OFN98_n232), 
	.B1(n565), 
	.B0(n47), 
	.A1(new_sboxw[19]), 
	.A0(n11));
   XNOR2X1 U985 (.Y(n565), 
	.B(n1362), 
	.A(round_key[83]));
   OAI221XL U986 (.Y(n1253), 
	.C0(n593), 
	.B1(n465), 
	.B0(n1379), 
	.A1(n106), 
	.A0(n592));
   XNOR2X1 U987 (.Y(n592), 
	.B(block[79]), 
	.A(round_key[79]));
   AOI222X1 U988 (.Y(n593), 
	.C1(n595), 
	.C0(FE_OFN97_n232), 
	.B1(n594), 
	.B0(n49), 
	.A1(new_sboxw[15]), 
	.A0(n11));
   XNOR2X1 U989 (.Y(n594), 
	.B(n1368), 
	.A(round_key[79]));
   OAI221XL U990 (.Y(n1248), 
	.C0(n556), 
	.B1(n465), 
	.B0(n1363), 
	.A1(n106), 
	.A0(n555));
   XNOR2X1 U991 (.Y(n555), 
	.B(block[84]), 
	.A(round_key[84]));
   AOI222X1 U992 (.Y(n556), 
	.C1(n558), 
	.C0(FE_OFN97_n232), 
	.B1(n557), 
	.B0(n46), 
	.A1(new_sboxw[20]), 
	.A0(n11));
   XNOR2X1 U993 (.Y(n557), 
	.B(n1398), 
	.A(round_key[84]));
   OAI221XL U994 (.Y(n1316), 
	.C0(n1067), 
	.B1(n945), 
	.B0(n1423), 
	.A1(n107), 
	.A0(FE_PHN5101_n1066));
   XNOR2X1 U995 (.Y(n1066), 
	.B(block[16]), 
	.A(round_key[16]));
   AOI222X1 U996 (.Y(n1067), 
	.C1(n1069), 
	.C0(FE_OFN98_n232), 
	.B1(n1068), 
	.B0(n97), 
	.A1(new_sboxw[16]), 
	.A0(n8));
   XNOR2X1 U997 (.Y(n1068), 
	.B(n1421), 
	.A(round_key[16]));
   OAI221XL U998 (.Y(n1313), 
	.C0(n1044), 
	.B1(n945), 
	.B0(n1397), 
	.A1(n107), 
	.A0(FE_PHN5133_n1043));
   XNOR2X1 U999 (.Y(n1043), 
	.B(block[19]), 
	.A(round_key[19]));
   AOI222X1 U1000 (.Y(n1044), 
	.C1(n1046), 
	.C0(FE_OFN97_n232), 
	.B1(n1045), 
	.B0(n83), 
	.A1(new_sboxw[19]), 
	.A0(n8));
   XNOR2X1 U1001 (.Y(n1045), 
	.B(n1447), 
	.A(round_key[19]));
   OAI221XL U1002 (.Y(n1320), 
	.C0(n1091), 
	.B1(n945), 
	.B0(n1348), 
	.A1(n107), 
	.A0(FE_PHN5152_n1090));
   XNOR2X1 U1003 (.Y(n1090), 
	.B(block[12]), 
	.A(round_key[12]));
   AOI222X1 U1004 (.Y(n1091), 
	.C1(n1093), 
	.C0(FE_OFN97_n232), 
	.B1(n1092), 
	.B0(n97), 
	.A1(new_sboxw[12]), 
	.A0(n8));
   XNOR2X1 U1005 (.Y(n1092), 
	.B(n1365), 
	.A(round_key[12]));
   OAI221XL U1006 (.Y(n1218), 
	.C0(n332), 
	.B1(n230), 
	.B0(n1447), 
	.A1(n99), 
	.A0(n331));
   XNOR2X1 U1007 (.Y(n331), 
	.B(block[115]), 
	.A(round_key[115]));
   AOI222X1 U1008 (.Y(n332), 
	.C1(n334), 
	.C0(n232), 
	.B1(n333), 
	.B0(n96), 
	.A1(n13), 
	.A0(new_sboxw[19]));
   XNOR2X1 U1009 (.Y(n333), 
	.B(n1383), 
	.A(round_key[115]));
   OAI221XL U1010 (.Y(n1221), 
	.C0(n355), 
	.B1(n230), 
	.B0(n1421), 
	.A1(n105), 
	.A0(n354));
   XNOR2X1 U1011 (.Y(n354), 
	.B(block[112]), 
	.A(round_key[112]));
   AOI222X1 U1012 (.Y(n355), 
	.C1(n357), 
	.C0(FE_OFN98_n232), 
	.B1(n356), 
	.B0(n38), 
	.A1(n13), 
	.A0(new_sboxw[16]));
   XNOR2X1 U1013 (.Y(n356), 
	.B(n1427), 
	.A(round_key[112]));
   OAI221XL U1014 (.Y(n1292), 
	.C0(n880), 
	.B1(n706), 
	.B0(n1420), 
	.A1(n106), 
	.A0(n879));
   XNOR2X1 U1015 (.Y(n879), 
	.B(block[40]), 
	.A(round_key[40]));
   AOI222X1 U1016 (.Y(n880), 
	.C1(n882), 
	.C0(FE_OFN98_n232), 
	.B1(n881), 
	.B0(n97), 
	.A1(new_sboxw[8]), 
	.A0(n16));
   XNOR2X1 U1017 (.Y(n881), 
	.B(n1419), 
	.A(round_key[40]));
   OAI221XL U1018 (.Y(n1289), 
	.C0(n860), 
	.B1(n706), 
	.B0(n1345), 
	.A1(n107), 
	.A0(n859));
   XNOR2X1 U1019 (.Y(n859), 
	.B(block[43]), 
	.A(round_key[43]));
   AOI222X1 U1020 (.Y(n860), 
	.C1(n862), 
	.C0(FE_OFN98_n232), 
	.B1(n861), 
	.B0(n97), 
	.A1(new_sboxw[11]), 
	.A0(n16));
   XNOR2X1 U1021 (.Y(n861), 
	.B(n187), 
	.A(round_key[43]));
   OAI221XL U1022 (.Y(n1321), 
	.C0(n1099), 
	.B1(n945), 
	.B0(n1372), 
	.A1(n107), 
	.A0(FE_PHN5091_n1098));
   XNOR2X1 U1023 (.Y(n1098), 
	.B(block[11]), 
	.A(round_key[11]));
   AOI222X1 U1024 (.Y(n1099), 
	.C1(n1101), 
	.C0(FE_OFN97_n232), 
	.B1(FE_PHN5172_n1100), 
	.B0(n97), 
	.A1(new_sboxw[11]), 
	.A0(n7));
   XNOR2X1 U1025 (.Y(n1100), 
	.B(n1396), 
	.A(round_key[11]));
   OAI221XL U1026 (.Y(n1226), 
	.C0(n387), 
	.B1(n230), 
	.B0(n187), 
	.A1(n106), 
	.A0(n386));
   XNOR2X1 U1027 (.Y(n386), 
	.B(block[107]), 
	.A(round_key[107]));
   AOI222X1 U1028 (.Y(n387), 
	.C1(n389), 
	.C0(FE_OFN98_n232), 
	.B1(n388), 
	.B0(n38), 
	.A1(n12), 
	.A0(new_sboxw[11]));
   XNOR2X1 U1029 (.Y(n388), 
	.B(n1345), 
	.A(round_key[107]));
   OAI221XL U1030 (.Y(n1242), 
	.C0(n509), 
	.B1(n465), 
	.B0(n1440), 
	.A1(n464), 
	.A0(n141));
   AOI222X1 U1031 (.Y(n509), 
	.C1(n512), 
	.C0(round_key[90]), 
	.B1(n146), 
	.B0(n511), 
	.A1(n510), 
	.A0(FE_OFN98_n232));
   OAI2BB2X1 U1032 (.Y(n511), 
	.B1(FE_PHN157_n237), 
	.B0(n1440), 
	.A1N(block[90]), 
	.A0N(n113));
   OAI22X1 U1033 (.Y(n512), 
	.B1(n30), 
	.B0(new_block[90]), 
	.A1(n105), 
	.A0(block[90]));
   OAI221XL U1034 (.Y(n1243), 
	.C0(n517), 
	.B1(n465), 
	.B0(n1429), 
	.A1(n464), 
	.A0(n142));
   AOI222X1 U1035 (.Y(n517), 
	.C1(n520), 
	.C0(round_key[89]), 
	.B1(n134), 
	.B0(n519), 
	.A1(n518), 
	.A0(FE_OFN98_n232));
   OAI2BB2X1 U1036 (.Y(n519), 
	.B1(FE_PHN157_n237), 
	.B0(n1429), 
	.A1N(block[89]), 
	.A0N(n114));
   OAI22X1 U1037 (.Y(n520), 
	.B1(n30), 
	.B0(new_block[89]), 
	.A1(n105), 
	.A0(block[89]));
   OAI221XL U1038 (.Y(n1305), 
	.C0(n980), 
	.B1(n945), 
	.B0(n1448), 
	.A1(n3), 
	.A0(n144));
   AOI222X1 U1039 (.Y(n980), 
	.C1(n983), 
	.C0(round_key[27]), 
	.B1(n152), 
	.B0(n982), 
	.A1(n981), 
	.A0(FE_OFN97_n232));
   OAI2BB2X1 U1040 (.Y(n982), 
	.B1(FE_PHN157_n237), 
	.B0(n1448), 
	.A1N(block[27]), 
	.A0N(n113));
   OAI22X1 U1041 (.Y(n983), 
	.B1(FE_PHN157_n237), 
	.B0(new_block[27]), 
	.A1(n105), 
	.A0(block[27]));
   OAI221XL U1042 (.Y(n1284), 
	.C0(n828), 
	.B1(n706), 
	.B0(n1424), 
	.A1(n107), 
	.A0(n827));
   XNOR2X1 U1043 (.Y(n827), 
	.B(block[48]), 
	.A(round_key[48]));
   AOI222X1 U1044 (.Y(n828), 
	.C1(n830), 
	.C0(FE_OFN98_n232), 
	.B1(n829), 
	.B0(n97), 
	.A1(new_sboxw[16]), 
	.A0(n17));
   XNOR2X1 U1045 (.Y(n829), 
	.B(n1423), 
	.A(round_key[48]));
   OAI221XL U1046 (.Y(n1281), 
	.C0(n805), 
	.B1(n706), 
	.B0(n1362), 
	.A1(n236), 
	.A0(n804));
   XNOR2X1 U1047 (.Y(n804), 
	.B(block[51]), 
	.A(round_key[51]));
   AOI222X1 U1048 (.Y(n805), 
	.C1(n807), 
	.C0(FE_OFN98_n232), 
	.B1(n806), 
	.B0(n97), 
	.A1(new_sboxw[19]), 
	.A0(n17));
   XNOR2X1 U1049 (.Y(n806), 
	.B(n1397), 
	.A(round_key[51]));
   INVX1 U1050 (.Y(n175), 
	.A(FE_PHN114_sword_ctr_reg_1_));
   NOR2X1 U1051 (.Y(n943), 
	.B(sword_ctr_reg[0]), 
	.A(n175));
   NOR2X1 U1052 (.Y(n704), 
	.B(FE_PHN114_sword_ctr_reg_1_), 
	.A(n56));
   NOR2X1 U1053 (.Y(n1182), 
	.B(n56), 
	.A(n175));
   AOI22X1 U1054 (.Y(n208), 
	.B1(n15), 
	.B0(new_block[58]), 
	.A1(n9), 
	.A0(new_block[90]));
   AOI22X1 U1055 (.Y(n212), 
	.B1(n15), 
	.B0(new_block[54]), 
	.A1(n9), 
	.A0(new_block[86]));
   OAI221XL U1056 (.Y(sboxw[26]), 
	.C0(n208), 
	.B1(n1442), 
	.B0(n194), 
	.A1(n1444), 
	.A0(n193));
   AOI22X1 U1057 (.Y(n198), 
	.B1(n15), 
	.B0(new_block[38]), 
	.A1(n9), 
	.A0(FE_PHN309_Dout_70_));
   OAI221XL U1058 (.Y(sboxw[22]), 
	.C0(n212), 
	.B1(n1407), 
	.B0(n194), 
	.A1(n1408), 
	.A0(n193));
   OAI221XL U1059 (.Y(sboxw[6]), 
	.C0(n198), 
	.B1(n1354), 
	.B0(n194), 
	.A1(n944), 
	.A0(n193));
   INVX1 U1060 (.Y(n1364), 
	.A(new_block[100]));
   INVX1 U1061 (.Y(n1370), 
	.A(new_block[9]));
   INVX1 U1062 (.Y(n189), 
	.A(new_block[4]));
   INVX1 U1063 (.Y(n1419), 
	.A(new_block[104]));
   INVX1 U1064 (.Y(n1387), 
	.A(new_block[20]));
   INVX1 U1065 (.Y(n1385), 
	.A(new_block[116]));
   INVX1 U1066 (.Y(n1384), 
	.A(new_block[124]));
   INVX1 U1067 (.Y(n1346), 
	.A(new_block[108]));
   INVX1 U1068 (.Y(n1433), 
	.A(new_block[105]));
   INVX1 U1069 (.Y(n184), 
	.A(new_block[96]));
   INVX1 U1070 (.Y(n1386), 
	.A(new_block[28]));
   INVX1 U1071 (.Y(n1348), 
	.A(new_block[12]));
   INVX1 U1072 (.Y(n1421), 
	.A(new_block[112]));
   INVX1 U1073 (.Y(n1447), 
	.A(new_block[115]));
   AOI22X1 U1074 (.Y(n203), 
	.B1(n15), 
	.B0(new_block[62]), 
	.A1(n9), 
	.A0(new_block[94]));
   AOI22X1 U1075 (.Y(n221), 
	.B1(n14), 
	.B0(new_block[46]), 
	.A1(n173), 
	.A0(FE_PHN292_Dout_78_));
   OAI221XL U1076 (.Y(sboxw[30]), 
	.C0(n203), 
	.B1(n1406), 
	.B0(n194), 
	.A1(n1377), 
	.A0(n193));
   OAI221XL U1077 (.Y(sboxw[14]), 
	.C0(n221), 
	.B1(n229), 
	.B0(n194), 
	.A1(n1378), 
	.A0(n193));
   INVX1 U1078 (.Y(n1425), 
	.A(new_block[8]));
   INVX1 U1079 (.Y(n1343), 
	.A(new_block[97]));
   INVX1 U1080 (.Y(n1394), 
	.A(new_block[1]));
   INVX1 U1081 (.Y(n1351), 
	.A(new_block[101]));
   INVX1 U1082 (.Y(n190), 
	.A(new_block[109]));
   INVX1 U1083 (.Y(n1405), 
	.A(new_block[125]));
   INVX1 U1084 (.Y(n192), 
	.A(new_block[5]));
   INVX1 U1085 (.Y(n1382), 
	.A(new_block[99]));
   INVX1 U1086 (.Y(n1395), 
	.A(new_block[98]));
   INVX1 U1087 (.Y(n1454), 
	.A(new_block[2]));
   INVX1 U1088 (.Y(n1452), 
	.A(new_block[3]));
   INVX1 U1089 (.Y(n1342), 
	.A(new_block[0]));
   INVX1 U1090 (.Y(n1418), 
	.A(new_block[120]));
   INVX1 U1091 (.Y(n1376), 
	.A(new_block[29]));
   INVX1 U1092 (.Y(n1436), 
	.A(new_block[17]));
   INVX1 U1093 (.Y(n1402), 
	.A(new_block[21]));
   INVX1 U1094 (.Y(n1366), 
	.A(new_block[13]));
   INVX1 U1095 (.Y(n1432), 
	.A(new_block[113]));
   INVX1 U1096 (.Y(n1375), 
	.A(new_block[117]));
   INVX1 U1097 (.Y(n1455), 
	.A(new_block[10]));
   INVX1 U1098 (.Y(n1431), 
	.A(new_block[121]));
   INVX1 U1099 (.Y(n1361), 
	.A(new_block[106]));
   INVX1 U1100 (.Y(n1422), 
	.A(new_block[24]));
   INVX1 U1101 (.Y(n1435), 
	.A(new_block[25]));
   INVX1 U1102 (.Y(n1446), 
	.A(new_block[123]));
   INVX1 U1103 (.Y(n1445), 
	.A(new_block[18]));
   INVX1 U1104 (.Y(n1423), 
	.A(new_block[16]));
   INVX1 U1105 (.Y(n1397), 
	.A(new_block[19]));
   INVX1 U1106 (.Y(n1443), 
	.A(new_block[114]));
   INVX1 U1107 (.Y(n1372), 
	.A(new_block[11]));
   INVX1 U1108 (.Y(n187), 
	.A(new_block[107]));
   INVX1 U1109 (.Y(n1448), 
	.A(new_block[27]));
   AOI22X1 U1110 (.Y(n197), 
	.B1(n15), 
	.B0(new_block[39]), 
	.A1(n9), 
	.A0(new_block[71]));
   AOI22X1 U1111 (.Y(n202), 
	.B1(n15), 
	.B0(new_block[63]), 
	.A1(n9), 
	.A0(new_block[95]));
   AOI22X1 U1112 (.Y(n220), 
	.B1(n14), 
	.B0(FE_PHN3105_Dout_47_), 
	.A1(n173), 
	.A0(new_block[79]));
   AOI22X1 U1113 (.Y(n211), 
	.B1(n15), 
	.B0(new_block[55]), 
	.A1(n9), 
	.A0(new_block[87]));
   OAI221XL U1114 (.Y(sboxw[15]), 
	.C0(n220), 
	.B1(n1199), 
	.B0(n194), 
	.A1(n1368), 
	.A0(n193));
   OAI221XL U1115 (.Y(sboxw[23]), 
	.C0(n211), 
	.B1(n1415), 
	.B0(n194), 
	.A1(n1416), 
	.A0(n193));
   OAI221XL U1116 (.Y(sboxw[31]), 
	.C0(n202), 
	.B1(n1417), 
	.B0(n194), 
	.A1(n1380), 
	.A0(n193));
   OAI221XL U1117 (.Y(sboxw[7]), 
	.C0(n197), 
	.B1(n1357), 
	.B0(n194), 
	.A1(n1381), 
	.A0(n193));
   INVX1 U1118 (.Y(n1354), 
	.A(new_block[102]));
   INVX1 U1119 (.Y(n944), 
	.A(new_block[6]));
   INVX1 U1120 (.Y(n1408), 
	.A(new_block[22]));
   INVX1 U1121 (.Y(n1407), 
	.A(new_block[118]));
   INVX1 U1122 (.Y(n1442), 
	.A(new_block[122]));
   INVX1 U1123 (.Y(n1444), 
	.A(new_block[26]));
   INVX1 U1124 (.Y(n229), 
	.A(new_block[110]));
   INVX1 U1125 (.Y(n1406), 
	.A(new_block[126]));
   INVX1 U1126 (.Y(n1377), 
	.A(new_block[30]));
   INVX1 U1127 (.Y(n1378), 
	.A(new_block[14]));
   INVX1 U1128 (.Y(n1381), 
	.A(new_block[7]));
   INVX1 U1129 (.Y(n1415), 
	.A(new_block[119]));
   INVX1 U1130 (.Y(n1199), 
	.A(new_block[111]));
   INVX1 U1131 (.Y(n1417), 
	.A(new_block[127]));
   INVX1 U1132 (.Y(n1416), 
	.A(new_block[23]));
   INVX1 U1133 (.Y(n1380), 
	.A(new_block[31]));
   INVX1 U1134 (.Y(n1368), 
	.A(new_block[15]));
   INVX1 U1135 (.Y(n1357), 
	.A(new_block[103]));
   XOR2X1 U1136 (.Y(n581), 
	.B(n583), 
	.A(n582));
   XOR2X1 U1137 (.Y(n583), 
	.B(n523), 
	.A(n584));
   XNOR2X1 U1138 (.Y(n582), 
	.B(n585), 
	.A(new_block[89]));
   XNOR2X1 U1139 (.Y(n584), 
	.B(n473), 
	.A(new_block[48]));
   XOR2X1 U1140 (.Y(n676), 
	.B(n678), 
	.A(n677));
   XOR2X1 U1141 (.Y(n678), 
	.B(n539), 
	.A(n679));
   XNOR2X1 U1142 (.Y(n677), 
	.B(n680), 
	.A(new_block[90]));
   XNOR2X1 U1143 (.Y(n679), 
	.B(n496), 
	.A(new_block[11]));
   XOR2X1 U1144 (.Y(n932), 
	.B(n934), 
	.A(n933));
   XOR2X1 U1145 (.Y(n934), 
	.B(n780), 
	.A(n935));
   XNOR2X1 U1146 (.Y(n933), 
	.B(n936), 
	.A(new_block[56]));
   XNOR2X1 U1147 (.Y(n935), 
	.B(n757), 
	.A(new_block[105]));
   XOR2X1 U1148 (.Y(n917), 
	.B(n919), 
	.A(n918));
   XOR2X1 U1149 (.Y(n919), 
	.B(n780), 
	.A(n920));
   XNOR2X1 U1150 (.Y(n918), 
	.B(n921), 
	.A(new_block[58]));
   XNOR2X1 U1151 (.Y(n920), 
	.B(n737), 
	.A(new_block[107]));
   XOR2X1 U1152 (.Y(n1046), 
	.B(n1048), 
	.A(n1047));
   XOR2X1 U1153 (.Y(n1048), 
	.B(n986), 
	.A(n1049));
   XNOR2X1 U1154 (.Y(n1047), 
	.B(n1050), 
	.A(new_block[27]));
   XNOR2X1 U1155 (.Y(n1049), 
	.B(n953), 
	.A(new_block[114]));
   XOR2X1 U1156 (.Y(n1061), 
	.B(n1063), 
	.A(n1062));
   XOR2X1 U1157 (.Y(n1063), 
	.B(n1003), 
	.A(n1064));
   XNOR2X1 U1158 (.Y(n1062), 
	.B(n1065), 
	.A(new_block[25]));
   XNOR2X1 U1159 (.Y(n1064), 
	.B(n953), 
	.A(new_block[112]));
   XOR2X1 U1160 (.Y(n566), 
	.B(n568), 
	.A(n567));
   XOR2X1 U1161 (.Y(n568), 
	.B(n506), 
	.A(n569));
   XNOR2X1 U1162 (.Y(n567), 
	.B(n570), 
	.A(new_block[50]));
   XNOR2X1 U1163 (.Y(n569), 
	.B(n473), 
	.A(new_block[10]));
   XOR2X1 U1164 (.Y(n822), 
	.B(n824), 
	.A(n823));
   XOR2X1 U1165 (.Y(n824), 
	.B(n764), 
	.A(n825));
   XNOR2X1 U1166 (.Y(n823), 
	.B(n826), 
	.A(new_block[16]));
   XNOR2X1 U1167 (.Y(n825), 
	.B(n714), 
	.A(new_block[104]));
   XOR2X1 U1168 (.Y(n807), 
	.B(n809), 
	.A(n808));
   XOR2X1 U1169 (.Y(n809), 
	.B(n747), 
	.A(n810));
   XNOR2X1 U1170 (.Y(n808), 
	.B(n811), 
	.A(new_block[18]));
   XNOR2X1 U1171 (.Y(n810), 
	.B(n714), 
	.A(new_block[106]));
   XOR2X1 U1172 (.Y(n691), 
	.B(n693), 
	.A(n692));
   XOR2X1 U1173 (.Y(n693), 
	.B(n539), 
	.A(n694));
   XNOR2X1 U1174 (.Y(n692), 
	.B(n695), 
	.A(new_block[96]));
   XNOR2X1 U1175 (.Y(n694), 
	.B(n516), 
	.A(new_block[88]));
   XOR2X1 U1176 (.Y(n1156), 
	.B(n1158), 
	.A(n1157));
   XOR2X1 U1177 (.Y(n1158), 
	.B(n1019), 
	.A(n1159));
   XNOR2X1 U1178 (.Y(n1157), 
	.B(n1160), 
	.A(new_block[34]));
   XNOR2X1 U1179 (.Y(n1159), 
	.B(n976), 
	.A(new_block[26]));
   XOR2X1 U1180 (.Y(n1171), 
	.B(n1173), 
	.A(n1172));
   XOR2X1 U1181 (.Y(n1173), 
	.B(n1019), 
	.A(n1174));
   XNOR2X1 U1182 (.Y(n1172), 
	.B(n1175), 
	.A(new_block[32]));
   XNOR2X1 U1183 (.Y(n1174), 
	.B(n996), 
	.A(new_block[24]));
   XOR2X1 U1184 (.Y(n467), 
	.B(n471), 
	.A(n470));
   XOR2X1 U1185 (.Y(n471), 
	.B(n473), 
	.A(n472));
   XNOR2X1 U1186 (.Y(n470), 
	.B(new_block[103]), 
	.A(n170));
   XOR2X1 U1187 (.Y(n742), 
	.B(n746), 
	.A(n745));
   XOR2X1 U1188 (.Y(n746), 
	.B(n748), 
	.A(n747));
   XOR2X1 U1189 (.Y(n745), 
	.B(n749), 
	.A(n738));
   XNOR2X1 U1190 (.Y(n749), 
	.B(new_block[19]), 
	.A(n151));
   XOR2X1 U1191 (.Y(n501), 
	.B(n505), 
	.A(n504));
   XOR2X1 U1192 (.Y(n505), 
	.B(n507), 
	.A(n506));
   XOR2X1 U1193 (.Y(n504), 
	.B(n508), 
	.A(n497));
   XNOR2X1 U1194 (.Y(n508), 
	.B(new_block[51]), 
	.A(n150));
   XOR2X1 U1195 (.Y(n981), 
	.B(n985), 
	.A(n984));
   XOR2X1 U1196 (.Y(n985), 
	.B(n987), 
	.A(n986));
   XOR2X1 U1197 (.Y(n984), 
	.B(n988), 
	.A(n977));
   XNOR2X1 U1198 (.Y(n988), 
	.B(new_block[115]), 
	.A(n152));
   XOR2X1 U1199 (.Y(n269), 
	.B(n273), 
	.A(n272));
   XOR2X1 U1200 (.Y(n273), 
	.B(n275), 
	.A(n274));
   XOR2X1 U1201 (.Y(n272), 
	.B(n276), 
	.A(n265));
   XNOR2X1 U1202 (.Y(n276), 
	.B(new_block[83]), 
	.A(n149));
   XOR2X1 U1203 (.Y(n990), 
	.B(n994), 
	.A(n993));
   XOR2X1 U1204 (.Y(n994), 
	.B(n996), 
	.A(n995));
   XNOR2X1 U1205 (.Y(n993), 
	.B(new_block[114]), 
	.A(n148));
   XOR2X1 U1206 (.Y(n278), 
	.B(n282), 
	.A(n281));
   XOR2X1 U1207 (.Y(n282), 
	.B(n284), 
	.A(n283));
   XNOR2X1 U1208 (.Y(n281), 
	.B(new_block[82]), 
	.A(n145));
   XOR2X1 U1209 (.Y(n510), 
	.B(n514), 
	.A(n513));
   XOR2X1 U1210 (.Y(n514), 
	.B(n516), 
	.A(n515));
   XNOR2X1 U1211 (.Y(n513), 
	.B(new_block[50]), 
	.A(n146));
   XOR2X1 U1212 (.Y(n751), 
	.B(n755), 
	.A(n754));
   XOR2X1 U1213 (.Y(n755), 
	.B(n757), 
	.A(n756));
   XNOR2X1 U1214 (.Y(n754), 
	.B(new_block[18]), 
	.A(n147));
   XOR2X1 U1215 (.Y(n759), 
	.B(n763), 
	.A(n762));
   XOR2X1 U1216 (.Y(n763), 
	.B(n765), 
	.A(n764));
   XOR2X1 U1217 (.Y(n762), 
	.B(n766), 
	.A(n738));
   XNOR2X1 U1218 (.Y(n766), 
	.B(new_block[17]), 
	.A(n135));
   XOR2X1 U1219 (.Y(n998), 
	.B(n1002), 
	.A(n1001));
   XOR2X1 U1220 (.Y(n1002), 
	.B(n1004), 
	.A(n1003));
   XOR2X1 U1221 (.Y(n1001), 
	.B(n1005), 
	.A(n977));
   XNOR2X1 U1222 (.Y(n1005), 
	.B(new_block[113]), 
	.A(n136));
   XOR2X1 U1223 (.Y(n286), 
	.B(n290), 
	.A(n289));
   XOR2X1 U1224 (.Y(n290), 
	.B(n292), 
	.A(n291));
   XOR2X1 U1225 (.Y(n289), 
	.B(n293), 
	.A(n265));
   XNOR2X1 U1226 (.Y(n293), 
	.B(new_block[81]), 
	.A(n133));
   XOR2X1 U1227 (.Y(n518), 
	.B(n522), 
	.A(n521));
   XOR2X1 U1228 (.Y(n522), 
	.B(n524), 
	.A(n523));
   XOR2X1 U1229 (.Y(n521), 
	.B(n525), 
	.A(n497));
   XNOR2X1 U1230 (.Y(n525), 
	.B(new_block[49]), 
	.A(n134));
   XOR2X1 U1231 (.Y(n527), 
	.B(n531), 
	.A(n530));
   XOR2X1 U1232 (.Y(n531), 
	.B(n532), 
	.A(n497));
   XNOR2X1 U1233 (.Y(n530), 
	.B(new_block[48]), 
	.A(n166));
   XOR2X1 U1234 (.Y(n1007), 
	.B(n1011), 
	.A(n1010));
   XOR2X1 U1235 (.Y(n1011), 
	.B(n1012), 
	.A(n977));
   XNOR2X1 U1236 (.Y(n1010), 
	.B(new_block[112]), 
	.A(n168));
   XOR2X1 U1237 (.Y(n295), 
	.B(n299), 
	.A(n298));
   XOR2X1 U1238 (.Y(n299), 
	.B(n300), 
	.A(n265));
   XNOR2X1 U1239 (.Y(n298), 
	.B(new_block[80]), 
	.A(n165));
   XOR2X1 U1240 (.Y(n233), 
	.B(n239), 
	.A(n238));
   XOR2X1 U1241 (.Y(n239), 
	.B(n241), 
	.A(n240));
   XNOR2X1 U1242 (.Y(n238), 
	.B(new_block[7]), 
	.A(n169));
   XOR2X1 U1243 (.Y(n475), 
	.B(n479), 
	.A(n478));
   XOR2X1 U1244 (.Y(n479), 
	.B(n481), 
	.A(n480));
   XNOR2X1 U1245 (.Y(n478), 
	.B(new_block[54]), 
	.A(n162));
   XOR2X1 U1246 (.Y(n243), 
	.B(n247), 
	.A(n246));
   XOR2X1 U1247 (.Y(n247), 
	.B(n249), 
	.A(n248));
   XNOR2X1 U1248 (.Y(n246), 
	.B(new_block[86]), 
	.A(n161));
   XOR2X1 U1249 (.Y(n251), 
	.B(n255), 
	.A(n254));
   XOR2X1 U1250 (.Y(n255), 
	.B(n257), 
	.A(n256));
   XNOR2X1 U1251 (.Y(n254), 
	.B(new_block[85]), 
	.A(n157));
   XOR2X1 U1252 (.Y(n483), 
	.B(n487), 
	.A(n486));
   XOR2X1 U1253 (.Y(n487), 
	.B(n489), 
	.A(n488));
   XNOR2X1 U1254 (.Y(n486), 
	.B(new_block[53]), 
	.A(n158));
   XOR2X1 U1255 (.Y(n491), 
	.B(n495), 
	.A(n494));
   XOR2X1 U1256 (.Y(n495), 
	.B(n497), 
	.A(n496));
   XOR2X1 U1257 (.Y(n494), 
	.B(n499), 
	.A(n498));
   XNOR2X1 U1258 (.Y(n499), 
	.B(new_block[52]), 
	.A(n154));
   XOR2X1 U1259 (.Y(n768), 
	.B(n772), 
	.A(n771));
   XOR2X1 U1260 (.Y(n772), 
	.B(n773), 
	.A(n738));
   XNOR2X1 U1261 (.Y(n771), 
	.B(new_block[16]), 
	.A(n167));
   XOR2X1 U1262 (.Y(n708), 
	.B(n712), 
	.A(n711));
   XOR2X1 U1263 (.Y(n712), 
	.B(n714), 
	.A(n713));
   XNOR2X1 U1264 (.Y(n711), 
	.B(new_block[71]), 
	.A(n171));
   XOR2X1 U1265 (.Y(n716), 
	.B(n720), 
	.A(n719));
   XOR2X1 U1266 (.Y(n720), 
	.B(n722), 
	.A(n721));
   XNOR2X1 U1267 (.Y(n719), 
	.B(new_block[22]), 
	.A(n163));
   XOR2X1 U1268 (.Y(n724), 
	.B(n728), 
	.A(n727));
   XOR2X1 U1269 (.Y(n728), 
	.B(n730), 
	.A(n729));
   XNOR2X1 U1270 (.Y(n727), 
	.B(new_block[21]), 
	.A(n159));
   XOR2X1 U1271 (.Y(n732), 
	.B(n736), 
	.A(n735));
   XOR2X1 U1272 (.Y(n736), 
	.B(n738), 
	.A(n737));
   XOR2X1 U1273 (.Y(n735), 
	.B(n740), 
	.A(n739));
   XNOR2X1 U1274 (.Y(n740), 
	.B(new_block[20]), 
	.A(n155));
   XOR2X1 U1275 (.Y(n971), 
	.B(n975), 
	.A(n974));
   XOR2X1 U1276 (.Y(n975), 
	.B(n977), 
	.A(n976));
   XOR2X1 U1277 (.Y(n974), 
	.B(n979), 
	.A(n978));
   XNOR2X1 U1278 (.Y(n979), 
	.B(new_block[116]), 
	.A(n156));
   XOR2X1 U1279 (.Y(n259), 
	.B(n263), 
	.A(n262));
   XOR2X1 U1280 (.Y(n263), 
	.B(n265), 
	.A(n264));
   XOR2X1 U1281 (.Y(n262), 
	.B(n267), 
	.A(n266));
   XNOR2X1 U1282 (.Y(n267), 
	.B(new_block[84]), 
	.A(n153));
   XOR2X1 U1283 (.Y(n947), 
	.B(n951), 
	.A(n950));
   XOR2X1 U1284 (.Y(n951), 
	.B(n953), 
	.A(n952));
   XNOR2X1 U1285 (.Y(n950), 
	.B(new_block[39]), 
	.A(n172));
   XOR2X1 U1286 (.Y(n955), 
	.B(n959), 
	.A(n958));
   XOR2X1 U1287 (.Y(n959), 
	.B(n961), 
	.A(n960));
   XNOR2X1 U1288 (.Y(n958), 
	.B(new_block[118]), 
	.A(n164));
   XOR2X1 U1289 (.Y(n963), 
	.B(n967), 
	.A(n966));
   XOR2X1 U1290 (.Y(n967), 
	.B(n969), 
	.A(n968));
   XNOR2X1 U1291 (.Y(n966), 
	.B(new_block[117]), 
	.A(n160));
   XOR2X1 U1292 (.Y(n334), 
	.B(n336), 
	.A(n335));
   XOR2X1 U1293 (.Y(n336), 
	.B(n274), 
	.A(n337));
   XNOR2X1 U1294 (.Y(n335), 
	.B(n338), 
	.A(new_block[42]));
   XNOR2X1 U1295 (.Y(n337), 
	.B(n241), 
	.A(new_block[123]));
   XOR2X1 U1296 (.Y(n349), 
	.B(n351), 
	.A(n350));
   XOR2X1 U1297 (.Y(n351), 
	.B(n291), 
	.A(n352));
   XNOR2X1 U1298 (.Y(n350), 
	.B(n353), 
	.A(new_block[40]));
   XNOR2X1 U1299 (.Y(n352), 
	.B(n241), 
	.A(new_block[121]));
   XOR2X1 U1300 (.Y(n799), 
	.B(n801), 
	.A(n800));
   XOR2X1 U1301 (.Y(n801), 
	.B(n739), 
	.A(n802));
   XNOR2X1 U1302 (.Y(n800), 
	.B(n803), 
	.A(new_block[19]));
   XNOR2X1 U1303 (.Y(n802), 
	.B(n714), 
	.A(new_block[107]));
   XOR2X1 U1304 (.Y(n1038), 
	.B(n1040), 
	.A(n1039));
   XOR2X1 U1305 (.Y(n1040), 
	.B(n978), 
	.A(n1041));
   XNOR2X1 U1306 (.Y(n1039), 
	.B(n1042), 
	.A(new_block[28]));
   XNOR2X1 U1307 (.Y(n1041), 
	.B(n953), 
	.A(new_block[115]));
   XOR2X1 U1308 (.Y(n326), 
	.B(n328), 
	.A(n327));
   XOR2X1 U1309 (.Y(n328), 
	.B(n266), 
	.A(n329));
   XNOR2X1 U1310 (.Y(n327), 
	.B(n330), 
	.A(new_block[43]));
   XNOR2X1 U1311 (.Y(n329), 
	.B(n241), 
	.A(new_block[124]));
   XOR2X1 U1312 (.Y(n444), 
	.B(n446), 
	.A(n445));
   XOR2X1 U1313 (.Y(n446), 
	.B(n307), 
	.A(n447));
   XNOR2X1 U1314 (.Y(n445), 
	.B(n448), 
	.A(new_block[2]));
   XNOR2X1 U1315 (.Y(n447), 
	.B(n264), 
	.A(new_block[122]));
   XOR2X1 U1316 (.Y(n436), 
	.B(n438), 
	.A(n437));
   XOR2X1 U1317 (.Y(n438), 
	.B(n307), 
	.A(n439));
   XNOR2X1 U1318 (.Y(n437), 
	.B(n440), 
	.A(new_block[3]));
   XNOR2X1 U1319 (.Y(n439), 
	.B(n257), 
	.A(new_block[123]));
   XOR2X1 U1320 (.Y(n558), 
	.B(n560), 
	.A(n559));
   XOR2X1 U1321 (.Y(n560), 
	.B(n498), 
	.A(n561));
   XNOR2X1 U1322 (.Y(n559), 
	.B(n562), 
	.A(new_block[51]));
   XNOR2X1 U1323 (.Y(n561), 
	.B(n473), 
	.A(new_block[11]));
   XOR2X1 U1324 (.Y(n668), 
	.B(n670), 
	.A(n669));
   XOR2X1 U1325 (.Y(n670), 
	.B(n539), 
	.A(n671));
   XNOR2X1 U1326 (.Y(n669), 
	.B(n672), 
	.A(new_block[91]));
   XNOR2X1 U1327 (.Y(n671), 
	.B(n489), 
	.A(new_block[12]));
   XOR2X1 U1328 (.Y(n909), 
	.B(n911), 
	.A(n910));
   XOR2X1 U1329 (.Y(n911), 
	.B(n780), 
	.A(n912));
   XNOR2X1 U1330 (.Y(n910), 
	.B(n913), 
	.A(new_block[59]));
   XNOR2X1 U1331 (.Y(n912), 
	.B(n730), 
	.A(new_block[108]));
   XOR2X1 U1332 (.Y(n459), 
	.B(n461), 
	.A(n460));
   XOR2X1 U1333 (.Y(n461), 
	.B(n307), 
	.A(n462));
   XNOR2X1 U1334 (.Y(n460), 
	.B(n463), 
	.A(new_block[120]));
   XNOR2X1 U1335 (.Y(n462), 
	.B(n284), 
	.A(new_block[0]));
   XOR2X1 U1336 (.Y(n1148), 
	.B(n1150), 
	.A(n1149));
   XOR2X1 U1337 (.Y(n1150), 
	.B(n1019), 
	.A(n1151));
   XNOR2X1 U1338 (.Y(n1149), 
	.B(n1152), 
	.A(new_block[35]));
   XNOR2X1 U1339 (.Y(n1151), 
	.B(n969), 
	.A(new_block[27]));
   XNOR2X1 U1340 (.Y(n780), 
	.B(new_block[71]), 
	.A(n1391));
   XNOR2X1 U1341 (.Y(n539), 
	.B(new_block[95]), 
	.A(n1357));
   XNOR2X1 U1342 (.Y(n307), 
	.B(new_block[7]), 
	.A(n1417));
   XNOR2X1 U1343 (.Y(n1019), 
	.B(new_block[39]), 
	.A(n1380));
   XNOR2X1 U1344 (.Y(n953), 
	.B(new_block[79]), 
	.A(n1415));
   XNOR2X1 U1345 (.Y(n241), 
	.B(new_block[87]), 
	.A(n1356));
   XNOR2X1 U1346 (.Y(n714), 
	.B(new_block[23]), 
	.A(n1199));
   XNOR2X1 U1347 (.Y(n473), 
	.B(new_block[55]), 
	.A(n1368));
   INVX1 U1348 (.Y(n705), 
	.A(new_block[38]));
   INVX1 U1349 (.Y(n1453), 
	.A(new_block[33]));
   INVX1 U1350 (.Y(n1374), 
	.A(new_block[44]));
   INVX1 U1351 (.Y(n191), 
	.A(new_block[37]));
   INVX1 U1352 (.Y(n1347), 
	.A(new_block[36]));
   XNOR2X1 U1353 (.Y(n857), 
	.B(new_block[71]), 
	.A(n1199));
   XNOR2X1 U1354 (.Y(n384), 
	.B(new_block[7]), 
	.A(n1356));
   XNOR2X1 U1355 (.Y(n1096), 
	.B(new_block[79]), 
	.A(n1341));
   XNOR2X1 U1356 (.Y(n616), 
	.B(new_block[15]), 
	.A(n1357));
   INVX1 U1357 (.Y(n1400), 
	.A(new_block[93]));
   INVX1 U1358 (.Y(n1399), 
	.A(new_block[92]));
   INVX1 U1359 (.Y(n1356), 
	.A(new_block[47]));
   INVX1 U1360 (.Y(n1353), 
	.A(new_block[46]));
   INVX1 U1361 (.Y(n1350), 
	.A(new_block[45]));
   OAI32X1 U1362 (.Y(n1336), 
	.B1(n182), 
	.B0(n1198), 
	.A2(n179), 
	.A1(FE_PHN2813_enc_round_nr_2_), 
	.A0(n181));
   INVX1 U1363 (.Y(n1371), 
	.A(new_block[74]));
   INVX1 U1364 (.Y(n185), 
	.A(new_block[65]));
   INVX1 U1365 (.Y(n1344), 
	.A(new_block[66]));
   INVX1 U1366 (.Y(n1369), 
	.A(new_block[72]));
   INVX1 U1367 (.Y(n1359), 
	.A(new_block[64]));
   INVX1 U1368 (.Y(n1396), 
	.A(new_block[75]));
   INVX1 U1369 (.Y(n1434), 
	.A(new_block[73]));
   INVX1 U1370 (.Y(n1401), 
	.A(new_block[77]));
   INVX1 U1371 (.Y(n1365), 
	.A(new_block[76]));
   INVX1 U1372 (.Y(n1349), 
	.A(new_block[68]));
   INVX1 U1373 (.Y(n1355), 
	.A(new_block[70]));
   INVX1 U1374 (.Y(n1352), 
	.A(new_block[69]));
   INVX1 U1375 (.Y(n1373), 
	.A(new_block[67]));
   INVX1 U1376 (.Y(n1410), 
	.A(new_block[94]));
   INVX1 U1377 (.Y(n1437), 
	.A(new_block[57]));
   INVX1 U1378 (.Y(n1390), 
	.A(new_block[62]));
   INVX1 U1379 (.Y(n1389), 
	.A(new_block[61]));
   INVX1 U1380 (.Y(n1388), 
	.A(new_block[60]));
   INVX1 U1381 (.Y(n1367), 
	.A(new_block[78]));
   INVX1 U1382 (.Y(n1360), 
	.A(new_block[41]));
   INVX1 U1383 (.Y(n1413), 
	.A(new_block[55]));
   INVX1 U1384 (.Y(n1409), 
	.A(new_block[54]));
   INVX1 U1385 (.Y(n1393), 
	.A(new_block[32]));
   INVX1 U1386 (.Y(n1451), 
	.A(new_block[34]));
   INVX1 U1387 (.Y(n188), 
	.A(new_block[35]));
   INVX1 U1388 (.Y(n1391), 
	.A(new_block[63]));
   INVX1 U1389 (.Y(n1358), 
	.A(new_block[95]));
   INVX1 U1390 (.Y(n1428), 
	.A(new_block[49]));
   INVX1 U1391 (.Y(n1403), 
	.A(new_block[53]));
   INVX1 U1392 (.Y(n1398), 
	.A(new_block[52]));
   INVX1 U1393 (.Y(n1449), 
	.A(new_block[91]));
   INVX1 U1394 (.Y(n1426), 
	.A(new_block[88]));
   INVX1 U1395 (.Y(n1450), 
	.A(new_block[59]));
   INVX1 U1396 (.Y(n1438), 
	.A(new_block[58]));
   INVX1 U1397 (.Y(n1392), 
	.A(new_block[56]));
   XNOR2X1 U1398 (.Y(n497), 
	.B(new_block[95]), 
	.A(n1413));
   XNOR2X1 U1399 (.Y(n977), 
	.B(new_block[31]), 
	.A(n1415));
   XNOR2X1 U1400 (.Y(n265), 
	.B(new_block[87]), 
	.A(n1417));
   XNOR2X1 U1401 (.Y(n738), 
	.B(new_block[63]), 
	.A(n1416));
   INVX1 U1402 (.Y(n1383), 
	.A(new_block[83]));
   INVX1 U1403 (.Y(n1441), 
	.A(new_block[82]));
   INVX1 U1404 (.Y(n1430), 
	.A(new_block[81]));
   INVX1 U1405 (.Y(n1427), 
	.A(new_block[80]));
   INVX1 U1406 (.Y(n1411), 
	.A(new_block[86]));
   INVX1 U1407 (.Y(n1363), 
	.A(new_block[84]));
   INVX1 U1408 (.Y(n1404), 
	.A(new_block[85]));
   INVX1 U1409 (.Y(n1379), 
	.A(new_block[79]));
   INVX1 U1410 (.Y(n186), 
	.A(new_block[42]));
   INVX1 U1411 (.Y(n1345), 
	.A(new_block[43]));
   INVX1 U1412 (.Y(n1440), 
	.A(new_block[90]));
   INVX1 U1413 (.Y(n1429), 
	.A(new_block[89]));
   INVX1 U1414 (.Y(n1341), 
	.A(new_block[39]));
   INVX1 U1415 (.Y(n1439), 
	.A(new_block[50]));
   INVX1 U1416 (.Y(n1424), 
	.A(new_block[48]));
   INVX1 U1417 (.Y(n1362), 
	.A(new_block[51]));
   NAND3X1 U1418 (.Y(n1194), 
	.C(next), 
	.B(n178), 
	.A(n180));
   OAI21XL U1419 (.Y(n1200), 
	.B0(n1201), 
	.A1(n180), 
	.A0(round[0]));
   NOR2X1 U1420 (.Y(n1197), 
	.B(n180), 
	.A(n54));
   XNOR2X1 U1421 (.Y(n532), 
	.B(new_block[96]), 
	.A(n1425));
   XNOR2X1 U1422 (.Y(n523), 
	.B(new_block[9]), 
	.A(n1343));
   XNOR2X1 U1423 (.Y(n498), 
	.B(new_block[12]), 
	.A(n1364));
   XNOR2X1 U1424 (.Y(n291), 
	.B(new_block[41]), 
	.A(n1394));
   XNOR2X1 U1425 (.Y(n516), 
	.B(new_block[89]), 
	.A(n1428));
   XNOR2X1 U1426 (.Y(n507), 
	.B(new_block[90]), 
	.A(n1439));
   XNOR2X1 U1427 (.Y(n748), 
	.B(new_block[58]), 
	.A(n1445));
   XNOR2X1 U1428 (.Y(n488), 
	.B(new_block[13]), 
	.A(n1351));
   XNOR2X1 U1429 (.Y(n300), 
	.B(new_block[40]), 
	.A(n1342));
   XNOR2X1 U1430 (.Y(n729), 
	.B(new_block[69]), 
	.A(n190));
   XNOR2X1 U1431 (.Y(n284), 
	.B(new_block[81]), 
	.A(n1431));
   XNOR2X1 U1432 (.Y(n257), 
	.B(new_block[84]), 
	.A(n1384));
   XNOR2X1 U1433 (.Y(n275), 
	.B(new_block[82]), 
	.A(n1442));
   XNOR2X1 U1434 (.Y(n249), 
	.B(new_block[85]), 
	.A(n1405));
   XNOR2X1 U1435 (.Y(n757), 
	.B(new_block[57]), 
	.A(n1436));
   XNOR2X1 U1436 (.Y(n730), 
	.B(new_block[60]), 
	.A(n1387));
   XNOR2X1 U1437 (.Y(n489), 
	.B(new_block[92]), 
	.A(n1398));
   XNOR2X1 U1438 (.Y(n481), 
	.B(new_block[93]), 
	.A(n1403));
   XNOR2X1 U1439 (.Y(n722), 
	.B(new_block[61]), 
	.A(n1402));
   XNOR2X1 U1440 (.Y(n987), 
	.B(new_block[26]), 
	.A(n1443));
   XNOR2X1 U1441 (.Y(n996), 
	.B(new_block[25]), 
	.A(n1432));
   XNOR2X1 U1442 (.Y(n969), 
	.B(new_block[28]), 
	.A(n1385));
   XNOR2X1 U1443 (.Y(n1003), 
	.B(new_block[73]), 
	.A(n1453));
   XNOR2X1 U1444 (.Y(n978), 
	.B(new_block[76]), 
	.A(n1347));
   XNOR2X1 U1445 (.Y(n266), 
	.B(new_block[4]), 
	.A(n1374));
   XNOR2X1 U1446 (.Y(n773), 
	.B(new_block[64]), 
	.A(n1419));
   XNOR2X1 U1447 (.Y(n1012), 
	.B(new_block[72]), 
	.A(n1393));
   XNOR2X1 U1448 (.Y(n739), 
	.B(new_block[68]), 
	.A(n1346));
   XNOR2X1 U1449 (.Y(n764), 
	.B(new_block[65]), 
	.A(n1433));
   XNOR2X1 U1450 (.Y(n968), 
	.B(new_block[77]), 
	.A(n191));
   XNOR2X1 U1451 (.Y(n256), 
	.B(new_block[5]), 
	.A(n1350));
   XNOR2X1 U1452 (.Y(n961), 
	.B(new_block[29]), 
	.A(n1375));
   XNOR2X1 U1453 (.Y(n765), 
	.B(new_block[56]), 
	.A(n1423));
   XNOR2X1 U1454 (.Y(n524), 
	.B(new_block[88]), 
	.A(n1424));
   XNOR2X1 U1455 (.Y(n496), 
	.B(new_block[91]), 
	.A(n1362));
   XNOR2X1 U1456 (.Y(n737), 
	.B(new_block[59]), 
	.A(n1397));
   XNOR2X1 U1457 (.Y(n976), 
	.B(new_block[27]), 
	.A(n1447));
   XNOR2X1 U1458 (.Y(n480), 
	.B(new_block[14]), 
	.A(n1354));
   XNOR2X1 U1459 (.Y(n292), 
	.B(new_block[80]), 
	.A(n1418));
   XNOR2X1 U1460 (.Y(n721), 
	.B(new_block[70]), 
	.A(n229));
   XNOR2X1 U1461 (.Y(n274), 
	.B(new_block[43]), 
	.A(n1452));
   XNOR2X1 U1462 (.Y(n1004), 
	.B(new_block[24]), 
	.A(n1421));
   XNOR2X1 U1463 (.Y(n264), 
	.B(new_block[83]), 
	.A(n1446));
   XNOR2X1 U1464 (.Y(n240), 
	.B(new_block[86]), 
	.A(n1406));
   XNOR2X1 U1465 (.Y(n960), 
	.B(new_block[78]), 
	.A(n705));
   XNOR2X1 U1466 (.Y(n472), 
	.B(new_block[94]), 
	.A(n1409));
   XNOR2X1 U1467 (.Y(n713), 
	.B(new_block[62]), 
	.A(n1408));
   XNOR2X1 U1468 (.Y(n283), 
	.B(new_block[42]), 
	.A(n1454));
   XNOR2X1 U1469 (.Y(n986), 
	.B(new_block[75]), 
	.A(n188));
   XNOR2X1 U1470 (.Y(n506), 
	.B(new_block[99]), 
	.A(n1372));
   XNOR2X1 U1471 (.Y(n747), 
	.B(new_block[67]), 
	.A(n187));
   XNOR2X1 U1472 (.Y(n515), 
	.B(new_block[98]), 
	.A(n1455));
   XNOR2X1 U1473 (.Y(n248), 
	.B(new_block[6]), 
	.A(n1353));
   XNOR2X1 U1474 (.Y(n995), 
	.B(new_block[74]), 
	.A(n1451));
   XNOR2X1 U1475 (.Y(n756), 
	.B(new_block[66]), 
	.A(n1361));
   XNOR2X1 U1476 (.Y(n952), 
	.B(new_block[30]), 
	.A(n1407));
   AOI21X1 U1477 (.Y(n1198), 
	.B0(n1200), 
	.A1(FE_PHN3408_enc_ctrl_reg_0_), 
	.A0(n181));
   OAI2BB2X1 U1478 (.Y(n1337), 
	.B1(n179), 
	.B0(round[1]), 
	.A1N(round[1]), 
	.A0N(n1200));
   OAI2BB1X1 U1479 (.Y(n1335), 
	.B0(n1196), 
	.A1N(round[3]), 
	.A0N(n1195));
   NAND4XL U1480 (.Y(n1196), 
	.D(n183), 
	.C(FE_PHN602_n1197), 
	.B(round[1]), 
	.A(FE_PHN2813_enc_round_nr_2_));
   OAI21XL U1481 (.Y(n1195), 
	.B0(n1198), 
	.A1(FE_PHN2813_enc_round_nr_2_), 
	.A0(n180));
   OAI2BB1X1 U1482 (.Y(n1334), 
	.B0(FE_PHN157_n237), 
	.A1N(n1194), 
	.A0N(ready));
   INVX1 U1483 (.Y(n1414), 
	.A(new_block[87]));
   INVX1 U1484 (.Y(n1420), 
	.A(new_block[40]));
   INVX1 U1485 (.Y(n1412), 
	.A(new_block[71]));
   OAI2BB1X1 U1486 (.Y(enc_ctrl_we), 
	.B0(n1205), 
	.A1N(n1193), 
	.A0N(n1182));
   OAI22X1 U1487 (.Y(n1205), 
	.B1(FE_PHN3408_enc_ctrl_reg_0_), 
	.B0(next), 
	.A1(FE_PHN3408_enc_ctrl_reg_0_), 
	.A0(n178));
endmodule

module aes_key_mem (
	clk, 
	reset_n, 
	key, 
	init, 
	round, 
	round_key, 
	ready, 
	sboxw, 
	new_sboxw, 
	FE_OFN37_reset_n, 
	FE_OFN39_reset_n, 
	FE_OFN40_reset_n, 
	FE_OFN42_reset_n, 
	FE_OFN43_reset_n, 
	FE_OFN44_reset_n, 
	FE_OFN45_reset_n, 
	FE_OFN46_reset_n, 
	FE_OFN47_reset_n, 
	FE_OFN48_reset_n, 
	FE_OFN53_reset_n, 
	FE_OFN55_reset_n, 
	FE_OFN58_reset_n, 
	clk_48Mhz__L6_N1, 
	clk_48Mhz__L6_N10, 
	clk_48Mhz__L6_N11, 
	clk_48Mhz__L6_N12, 
	clk_48Mhz__L6_N13, 
	clk_48Mhz__L6_N14, 
	clk_48Mhz__L6_N15, 
	clk_48Mhz__L6_N16, 
	clk_48Mhz__L6_N17, 
	clk_48Mhz__L6_N18, 
	clk_48Mhz__L6_N19, 
	clk_48Mhz__L6_N2, 
	clk_48Mhz__L6_N20, 
	clk_48Mhz__L6_N21, 
	clk_48Mhz__L6_N22, 
	clk_48Mhz__L6_N23, 
	clk_48Mhz__L6_N24, 
	clk_48Mhz__L6_N25, 
	clk_48Mhz__L6_N26, 
	clk_48Mhz__L6_N27, 
	clk_48Mhz__L6_N28, 
	clk_48Mhz__L6_N29, 
	clk_48Mhz__L6_N3, 
	clk_48Mhz__L6_N30, 
	clk_48Mhz__L6_N31, 
	clk_48Mhz__L6_N32, 
	clk_48Mhz__L6_N33, 
	clk_48Mhz__L6_N34, 
	clk_48Mhz__L6_N35, 
	clk_48Mhz__L6_N36, 
	clk_48Mhz__L6_N37, 
	clk_48Mhz__L6_N38, 
	clk_48Mhz__L6_N4, 
	clk_48Mhz__L6_N42, 
	clk_48Mhz__L6_N43, 
	clk_48Mhz__L6_N44, 
	clk_48Mhz__L6_N45, 
	clk_48Mhz__L6_N46, 
	clk_48Mhz__L6_N47, 
	clk_48Mhz__L6_N5, 
	clk_48Mhz__L6_N6, 
	clk_48Mhz__L6_N7, 
	clk_48Mhz__L6_N8, 
	clk_48Mhz__L6_N9);
   input clk;
   input reset_n;
   input [127:0] key;
   input init;
   input [3:0] round;
   output [127:0] round_key;
   output ready;
   output [31:0] sboxw;
   input [31:0] new_sboxw;
   input FE_OFN37_reset_n;
   input FE_OFN39_reset_n;
   input FE_OFN40_reset_n;
   input FE_OFN42_reset_n;
   input FE_OFN43_reset_n;
   input FE_OFN44_reset_n;
   input FE_OFN45_reset_n;
   input FE_OFN46_reset_n;
   input FE_OFN47_reset_n;
   input FE_OFN48_reset_n;
   input FE_OFN53_reset_n;
   input FE_OFN55_reset_n;
   input FE_OFN58_reset_n;
   input clk_48Mhz__L6_N1;
   input clk_48Mhz__L6_N10;
   input clk_48Mhz__L6_N11;
   input clk_48Mhz__L6_N12;
   input clk_48Mhz__L6_N13;
   input clk_48Mhz__L6_N14;
   input clk_48Mhz__L6_N15;
   input clk_48Mhz__L6_N16;
   input clk_48Mhz__L6_N17;
   input clk_48Mhz__L6_N18;
   input clk_48Mhz__L6_N19;
   input clk_48Mhz__L6_N2;
   input clk_48Mhz__L6_N20;
   input clk_48Mhz__L6_N21;
   input clk_48Mhz__L6_N22;
   input clk_48Mhz__L6_N23;
   input clk_48Mhz__L6_N24;
   input clk_48Mhz__L6_N25;
   input clk_48Mhz__L6_N26;
   input clk_48Mhz__L6_N27;
   input clk_48Mhz__L6_N28;
   input clk_48Mhz__L6_N29;
   input clk_48Mhz__L6_N3;
   input clk_48Mhz__L6_N30;
   input clk_48Mhz__L6_N31;
   input clk_48Mhz__L6_N32;
   input clk_48Mhz__L6_N33;
   input clk_48Mhz__L6_N34;
   input clk_48Mhz__L6_N35;
   input clk_48Mhz__L6_N36;
   input clk_48Mhz__L6_N37;
   input clk_48Mhz__L6_N38;
   input clk_48Mhz__L6_N4;
   input clk_48Mhz__L6_N42;
   input clk_48Mhz__L6_N43;
   input clk_48Mhz__L6_N44;
   input clk_48Mhz__L6_N45;
   input clk_48Mhz__L6_N46;
   input clk_48Mhz__L6_N47;
   input clk_48Mhz__L6_N5;
   input clk_48Mhz__L6_N6;
   input clk_48Mhz__L6_N7;
   input clk_48Mhz__L6_N8;
   input clk_48Mhz__L6_N9;

   // Internal wires
   wire FE_PHN5077_n2415;
   wire FE_PHN5076_n2407;
   wire FE_PHN5073_n2430;
   wire FE_PHN5066_n2407;
   wire FE_PHN5065_n2415;
   wire FE_PHN5063_n2400;
   wire FE_PHN5062_n2416;
   wire FE_PHN5061_n2391;
   wire FE_PHN5060_n2408;
   wire FE_PHN5058_n2392;
   wire FE_PHN5057_n2399;
   wire FE_PHN5056_n2412;
   wire FE_PHN5055_n2409;
   wire FE_PHN5054_n2403;
   wire FE_PHN5053_n2393;
   wire FE_PHN5052_n2417;
   wire FE_PHN5051_n2404;
   wire FE_PHN5050_n2411;
   wire FE_PHN5049_n2401;
   wire FE_PHN5047_n2431;
   wire FE_PHN5044_n2397;
   wire FE_PHN5043_n2406;
   wire FE_PHN5042_n2394;
   wire FE_PHN5041_n2398;
   wire FE_PHN5040_n2410;
   wire FE_PHN5039_n2405;
   wire FE_PHN5038_n2420;
   wire FE_PHN5037_n2402;
   wire FE_PHN5036_n2359;
   wire FE_PHN5035_n2419;
   wire FE_PHN5034_n2351;
   wire FE_PHN5033_n2414;
   wire FE_PHN5032_n2390;
   wire FE_PHN5031_n2413;
   wire FE_PHN5030_n2418;
   wire FE_PHN5029_n2352;
   wire FE_PHN5028_n2363;
   wire FE_PHN5027_n2396;
   wire FE_PHN5026_n2353;
   wire FE_PHN5025_n2354;
   wire FE_PHN5024_n2344;
   wire FE_PHN5023_n2293;
   wire FE_PHN5022_n2356;
   wire FE_PHN5021_n2297;
   wire FE_PHN5020_n2395;
   wire FE_PHN5019_n2349;
   wire FE_PHN5018_n2300;
   wire FE_PHN5017_n2362;
   wire FE_PHN5016_n2335;
   wire FE_PHN5015_n2360;
   wire FE_PHN5014_n2295;
   wire FE_PHN5013_n2346;
   wire FE_PHN5012_n2345;
   wire FE_PHN5011_n2336;
   wire FE_PHN5010_n2357;
   wire FE_PHN5009_n2361;
   wire FE_PHN5008_n2348;
   wire FE_PHN5007_n2341;
   wire FE_PHN5006_n2364;
   wire FE_PHN5005_n2296;
   wire FE_PHN5004_n2339;
   wire FE_PHN5003_n2340;
   wire FE_PHN5002_n2347;
   wire FE_PHN5001_n2342;
   wire FE_PHN5000_n2343;
   wire FE_PHN4999_n2338;
   wire FE_PHN4998_n2355;
   wire FE_PHN4997_n2389;
   wire FE_PHN4996_key_mem_846_;
   wire FE_PHN4995_n2334;
   wire FE_PHN4994_n2358;
   wire FE_PHN4993_n2294;
   wire FE_PHN4992_n2299;
   wire FE_PHN4991_n1210;
   wire FE_PHN4990_n2333;
   wire FE_PHN4989_n2337;
   wire FE_PHN4988_n1730;
   wire FE_PHN4987_n1916;
   wire FE_PHN4986_n2298;
   wire FE_PHN4985_n1981;
   wire FE_PHN4984_n2350;
   wire FE_PHN4983_n1052;
   wire FE_PHN4982_n1207;
   wire FE_PHN4981_n1178;
   wire FE_PHN4980_n2425;
   wire FE_PHN4979_n1085;
   wire FE_PHN4978_n1027;
   wire FE_PHN4977_n1329;
   wire FE_PHN4976_n1239;
   wire FE_PHN4975_n1246;
   wire FE_PHN4974_n1192;
   wire FE_PHN4973_n2304;
   wire FE_PHN4972_n1224;
   wire FE_PHN4971_n1020;
   wire FE_PHN4970_n957;
   wire FE_PHN4969_n1116;
   wire FE_PHN4968_n2312;
   wire FE_PHN4967_n1179;
   wire FE_PHN4966_n1067;
   wire FE_PHN4965_n918;
   wire FE_PHN4964_n1558;
   wire FE_PHN4963_n1073;
   wire FE_PHN4961_n1191;
   wire FE_PHN4960_n1118;
   wire FE_PHN4959_n1033;
   wire FE_PHN4958_n1062;
   wire FE_PHN4956_n1319;
   wire FE_PHN4955_n1390;
   wire FE_PHN4954_n2376;
   wire FE_PHN4953_n1978;
   wire FE_PHN4952_n931;
   wire FE_PHN4951_n1263;
   wire FE_PHN4950_n1612;
   wire FE_PHN4949_n1231;
   wire FE_PHN4948_n2379;
   wire FE_PHN4947_n1359;
   wire FE_PHN4946_n1208;
   wire FE_PHN4945_n1327;
   wire FE_PHN4944_n1268;
   wire FE_PHN4943_n1243;
   wire FE_PHN4942_n2385;
   wire FE_PHN4941_n1932;
   wire FE_PHN4940_n2370;
   wire FE_PHN4939_n965;
   wire FE_PHN4938_n992;
   wire FE_PHN4937_n1248;
   wire FE_PHN4936_n1308;
   wire FE_PHN4935_n1099;
   wire FE_PHN4934_n1173;
   wire FE_PHN4933_n1537;
   wire FE_PHN4932_n1126;
   wire FE_PHN4931_n981;
   wire FE_PHN4930_n1571;
   wire FE_PHN4929_n1233;
   wire FE_PHN4928_n2091;
   wire FE_PHN4927_n1621;
   wire FE_PHN4926_n1261;
   wire FE_PHN4925_n1038;
   wire FE_PHN4924_n1209;
   wire FE_PHN4923_n1154;
   wire FE_PHN4922_n1252;
   wire FE_PHN4921_n1267;
   wire FE_PHN4920_n1599;
   wire FE_PHN4919_n1152;
   wire FE_PHN4918_n1999;
   wire FE_PHN4917_n1247;
   wire FE_PHN4916_n1193;
   wire FE_PHN4915_n1180;
   wire FE_PHN4914_n1933;
   wire FE_PHN4913_n1048;
   wire FE_PHN4912_n1262;
   wire FE_PHN4911_n1253;
   wire FE_PHN4910_n1888;
   wire FE_PHN4909_n1149;
   wire FE_PHN4908_n1141;
   wire FE_PHN4907_n1256;
   wire FE_PHN4906_n1142;
   wire FE_PHN4905_n1607;
   wire FE_PHN4904_n1137;
   wire FE_PHN4903_n1194;
   wire FE_PHN4902_n1214;
   wire FE_PHN4901_n1886;
   wire FE_PHN4900_n1220;
   wire FE_PHN4899_n2365;
   wire FE_PHN4898_n1037;
   wire FE_PHN4897_n974;
   wire FE_PHN4896_n958;
   wire FE_PHN4895_n2428;
   wire FE_PHN4894_n1984;
   wire FE_PHN4893_n1186;
   wire FE_PHN4892_n1221;
   wire FE_PHN4891_n1198;
   wire FE_PHN4890_n1139;
   wire FE_PHN4889_n1086;
   wire FE_PHN4888_n2327;
   wire FE_PHN4887_n1371;
   wire FE_PHN4886_n1293;
   wire FE_PHN4885_n2229;
   wire FE_PHN4884_n2313;
   wire FE_PHN4883_n2017;
   wire FE_PHN4882_n1144;
   wire FE_PHN4881_n1586;
   wire FE_PHN4880_n1001;
   wire FE_PHN4879_n1232;
   wire FE_PHN4878_n1244;
   wire FE_PHN4877_n1965;
   wire FE_PHN4876_n2319;
   wire FE_PHN4875_n1989;
   wire FE_PHN4874_n2326;
   wire FE_PHN4873_n1021;
   wire FE_PHN4872_n1344;
   wire FE_PHN4871_n886;
   wire FE_PHN4870_n1045;
   wire FE_PHN4869_n1976;
   wire FE_PHN4868_n1563;
   wire FE_PHN4867_n1393;
   wire FE_PHN4866_n1943;
   wire FE_PHN4865_n1356;
   wire FE_PHN4864_n1598;
   wire FE_PHN4863_n1526;
   wire FE_PHN4862_n1106;
   wire FE_PHN4861_n1827;
   wire FE_PHN4860_n1087;
   wire FE_PHN4859_n935;
   wire FE_PHN4858_n1264;
   wire FE_PHN4857_n1304;
   wire FE_PHN4856_n1189;
   wire FE_PHN4855_n1230;
   wire FE_PHN4853_n1158;
   wire FE_PHN4852_n1649;
   wire FE_PHN4851_n2371;
   wire FE_PHN4850_n1203;
   wire FE_PHN4849_n2035;
   wire FE_PHN4848_n1165;
   wire FE_PHN4847_n1009;
   wire FE_PHN4846_n1115;
   wire FE_PHN4845_n2315;
   wire FE_PHN4844_n1647;
   wire FE_PHN4843_n1228;
   wire FE_PHN4842_n1251;
   wire FE_PHN4841_n1134;
   wire FE_PHN4840_n2332;
   wire FE_PHN4839_n1872;
   wire FE_PHN4838_n1282;
   wire FE_PHN4837_n1171;
   wire FE_PHN4836_n1501;
   wire FE_PHN4835_n2036;
   wire FE_PHN4834_n1070;
   wire FE_PHN4833_n1630;
   wire FE_PHN4832_n1617;
   wire FE_PHN4831_n1100;
   wire FE_PHN4830_n1614;
   wire FE_PHN4829_n1223;
   wire FE_PHN4828_n1608;
   wire FE_PHN4827_n954;
   wire FE_PHN4826_n1065;
   wire FE_PHN4825_n1632;
   wire FE_PHN4824_n1172;
   wire FE_PHN4823_n1204;
   wire FE_PHN4822_n1091;
   wire FE_PHN4821_n1962;
   wire FE_PHN4820_n1199;
   wire FE_PHN4819_n1148;
   wire FE_PHN4818_n1973;
   wire FE_PHN4817_n1348;
   wire FE_PHN4816_n1249;
   wire FE_PHN4815_n1156;
   wire FE_PHN4814_n2308;
   wire FE_PHN4813_n1355;
   wire FE_PHN4812_n2302;
   wire FE_PHN4811_n1241;
   wire FE_PHN4810_n1557;
   wire FE_PHN4809_n2366;
   wire FE_PHN4808_n1488;
   wire FE_PHN4807_n1681;
   wire FE_PHN4806_n1619;
   wire FE_PHN4805_n1300;
   wire FE_PHN4804_n1039;
   wire FE_PHN4803_n1587;
   wire FE_PHN4802_n1611;
   wire FE_PHN4801_n1307;
   wire FE_PHN4800_n1066;
   wire FE_PHN4799_n1326;
   wire FE_PHN4798_n969;
   wire FE_PHN4797_n1561;
   wire FE_PHN4796_n1206;
   wire FE_PHN4795_n2015;
   wire FE_PHN4794_n1636;
   wire FE_PHN4793_n1357;
   wire FE_PHN4792_n1643;
   wire FE_PHN4791_n1550;
   wire FE_PHN4790_n1237;
   wire FE_PHN4789_n1053;
   wire FE_PHN4788_n1912;
   wire FE_PHN4787_n2314;
   wire FE_PHN4786_n1922;
   wire FE_PHN4785_n1150;
   wire FE_PHN4784_n2022;
   wire FE_PHN4783_n2383;
   wire FE_PHN4782_n1164;
   wire FE_PHN4781_n1605;
   wire FE_PHN4780_n1294;
   wire FE_PHN4779_n1987;
   wire FE_PHN4778_n1043;
   wire FE_PHN4777_n1103;
   wire FE_PHN4776_n1651;
   wire FE_PHN4775_n902;
   wire FE_PHN4774_n1867;
   wire FE_PHN4773_n1980;
   wire FE_PHN4772_n1638;
   wire FE_PHN4771_n1529;
   wire FE_PHN4770_n1078;
   wire FE_PHN4769_n1129;
   wire FE_PHN4768_n1615;
   wire FE_PHN4767_n2369;
   wire FE_PHN4766_n1213;
   wire FE_PHN4765_n1157;
   wire FE_PHN4764_n1177;
   wire FE_PHN4763_n1302;
   wire FE_PHN4762_n1059;
   wire FE_PHN4761_n1276;
   wire FE_PHN4760_n1564;
   wire FE_PHN4759_n2024;
   wire FE_PHN4758_n1202;
   wire FE_PHN4757_n1216;
   wire FE_PHN4756_n926;
   wire FE_PHN4755_n1155;
   wire FE_PHN4754_n1584;
   wire FE_PHN4753_n1589;
   wire FE_PHN4752_n1019;
   wire FE_PHN4751_n920;
   wire FE_PHN4750_n1200;
   wire FE_PHN4749_n2114;
   wire FE_PHN4748_n1601;
   wire FE_PHN4747_n2004;
   wire FE_PHN4746_n1255;
   wire FE_PHN4745_n1979;
   wire FE_PHN4744_n1117;
   wire FE_PHN4743_n1349;
   wire FE_PHN4742_n1058;
   wire FE_PHN4741_n1940;
   wire FE_PHN4740_n1093;
   wire FE_PHN4739_n1354;
   wire FE_PHN4738_n1159;
   wire FE_PHN4737_n1642;
   wire FE_PHN4736_n1602;
   wire FE_PHN4735_n1629;
   wire FE_PHN4734_n2084;
   wire FE_PHN4733_n1215;
   wire FE_PHN4732_n973;
   wire FE_PHN4731_n2188;
   wire FE_PHN4730_n2180;
   wire FE_PHN4729_n1935;
   wire FE_PHN4728_n2033;
   wire FE_PHN4727_n1338;
   wire FE_PHN4726_n1195;
   wire FE_PHN4725_n1138;
   wire FE_PHN4724_n1365;
   wire FE_PHN4723_n1167;
   wire FE_PHN4722_n1990;
   wire FE_PHN4721_n1887;
   wire FE_PHN4720_n2256;
   wire FE_PHN4719_n1075;
   wire FE_PHN4718_n2209;
   wire FE_PHN4717_n1110;
   wire FE_PHN4716_n1622;
   wire FE_PHN4715_n2320;
   wire FE_PHN4714_n1284;
   wire FE_PHN4713_n1283;
   wire FE_PHN4712_n2031;
   wire FE_PHN4711_n1640;
   wire FE_PHN4710_n1131;
   wire FE_PHN4709_n915;
   wire FE_PHN4708_n1119;
   wire FE_PHN4707_n1205;
   wire FE_PHN4706_n1977;
   wire FE_PHN4705_n2117;
   wire FE_PHN4704_n1527;
   wire FE_PHN4703_n2375;
   wire FE_PHN4702_n1350;
   wire FE_PHN4701_n2424;
   wire FE_PHN4700_n1090;
   wire FE_PHN4699_n1147;
   wire FE_PHN4698_n1689;
   wire FE_PHN4697_n1585;
   wire FE_PHN4696_n953;
   wire FE_PHN4695_n1949;
   wire FE_PHN4694_n1125;
   wire FE_PHN4693_n1944;
   wire FE_PHN4692_n2201;
   wire FE_PHN4691_n1929;
   wire FE_PHN4690_n1641;
   wire FE_PHN4689_n2030;
   wire FE_PHN4688_n1551;
   wire FE_PHN4687_n1339;
   wire FE_PHN4686_n1183;
   wire FE_PHN4685_n1528;
   wire FE_PHN4684_n1746;
   wire FE_PHN4683_n2011;
   wire FE_PHN4682_n1392;
   wire FE_PHN4681_n1533;
   wire FE_PHN4680_n1130;
   wire FE_PHN4679_n1553;
   wire FE_PHN4678_n1303;
   wire FE_PHN4677_n1098;
   wire FE_PHN4676_n2060;
   wire FE_PHN4675_n1992;
   wire FE_PHN4674_n1315;
   wire FE_PHN4673_n2330;
   wire FE_PHN4672_n1235;
   wire FE_PHN4671_n925;
   wire FE_PHN4670_n1317;
   wire FE_PHN4669_n1419;
   wire FE_PHN4668_n1174;
   wire FE_PHN4667_n1212;
   wire FE_PHN4665_n2223;
   wire FE_PHN4664_n2324;
   wire FE_PHN4663_n1637;
   wire FE_PHN4662_n936;
   wire FE_PHN4661_n1324;
   wire FE_PHN4660_n1322;
   wire FE_PHN4659_n2016;
   wire FE_PHN4658_n2305;
   wire FE_PHN4657_n2116;
   wire FE_PHN4656_n1226;
   wire FE_PHN4655_n2081;
   wire FE_PHN4654_n1610;
   wire FE_PHN4653_n1069;
   wire FE_PHN4652_n1959;
   wire FE_PHN4651_n1566;
   wire FE_PHN4650_n2316;
   wire FE_PHN4649_n1108;
   wire FE_PHN4648_n1025;
   wire FE_PHN4647_n1036;
   wire FE_PHN4646_n1188;
   wire FE_PHN4644_n1532;
   wire FE_PHN4643_n1352;
   wire FE_PHN4642_n1569;
   wire FE_PHN4641_n1363;
   wire FE_PHN4640_n1120;
   wire FE_PHN4639_n1145;
   wire FE_PHN4638_n1123;
   wire FE_PHN4637_n1219;
   wire FE_PHN4636_n1321;
   wire FE_PHN4635_n1613;
   wire FE_PHN4634_n2119;
   wire FE_PHN4633_n1538;
   wire FE_PHN4632_n1915;
   wire FE_PHN4631_n2275;
   wire FE_PHN4630_n1575;
   wire FE_PHN4629_n2368;
   wire FE_PHN4628_n932;
   wire FE_PHN4627_n1072;
   wire FE_PHN4626_n1272;
   wire FE_PHN4625_n1570;
   wire FE_PHN4624_n1556;
   wire FE_PHN4623_n1836;
   wire FE_PHN4622_n1806;
   wire FE_PHN4621_n1924;
   wire FE_PHN4620_n1313;
   wire FE_PHN4619_n1026;
   wire FE_PHN4618_n1007;
   wire FE_PHN4617_n2014;
   wire FE_PHN4616_n2155;
   wire FE_PHN4615_n1281;
   wire FE_PHN4614_n907;
   wire FE_PHN4613_n1583;
   wire FE_PHN4612_n887;
   wire FE_PHN4611_n1525;
   wire FE_PHN4610_n1133;
   wire FE_PHN4609_n2019;
   wire FE_PHN4608_n2283;
   wire FE_PHN4607_n909;
   wire FE_PHN4606_n1381;
   wire FE_PHN4605_n1176;
   wire FE_PHN4604_n1136;
   wire FE_PHN4603_n2139;
   wire FE_PHN4602_n1548;
   wire FE_PHN4601_n1972;
   wire FE_PHN4600_n1182;
   wire FE_PHN4599_n1380;
   wire FE_PHN4598_n1582;
   wire FE_PHN4597_n960;
   wire FE_PHN4596_n977;
   wire FE_PHN4595_n1388;
   wire FE_PHN4594_n1934;
   wire FE_PHN4593_n1387;
   wire FE_PHN4592_n1543;
   wire FE_PHN4591_n2310;
   wire FE_PHN4590_n1332;
   wire FE_PHN4589_n948;
   wire FE_PHN4588_n2049;
   wire FE_PHN4587_n1744;
   wire FE_PHN4586_n1918;
   wire FE_PHN4585_n1970;
   wire FE_PHN4584_n1986;
   wire FE_PHN4583_n1211;
   wire FE_PHN4582_n1982;
   wire FE_PHN4581_n1623;
   wire FE_PHN4580_n1857;
   wire FE_PHN4579_n1018;
   wire FE_PHN4578_n1068;
   wire FE_PHN4577_n1812;
   wire FE_PHN4576_n1092;
   wire FE_PHN4575_n2309;
   wire FE_PHN4574_n1639;
   wire FE_PHN4573_n1015;
   wire FE_PHN4572_n2005;
   wire FE_PHN4571_n1914;
   wire FE_PHN4570_n2007;
   wire FE_PHN4569_n1132;
   wire FE_PHN4568_n1331;
   wire FE_PHN4567_n2185;
   wire FE_PHN4566_n1952;
   wire FE_PHN4565_n1820;
   wire FE_PHN4564_n2384;
   wire FE_PHN4563_n1966;
   wire FE_PHN4562_n2010;
   wire FE_PHN4561_n1044;
   wire FE_PHN4560_n1383;
   wire FE_PHN4559_n1190;
   wire FE_PHN4558_n1947;
   wire FE_PHN4557_n1181;
   wire FE_PHN4556_n1005;
   wire FE_PHN4555_n1245;
   wire FE_PHN4554_n999;
   wire FE_PHN4553_n1113;
   wire FE_PHN4552_n1360;
   wire FE_PHN4551_n1579;
   wire FE_PHN4550_n1559;
   wire FE_PHN4549_n1361;
   wire FE_PHN4548_n1534;
   wire FE_PHN4547_n2182;
   wire FE_PHN4546_n1080;
   wire FE_PHN4545_n1146;
   wire FE_PHN4544_n1004;
   wire FE_PHN4543_n1006;
   wire FE_PHN4542_n2046;
   wire FE_PHN4541_n1187;
   wire FE_PHN4540_n1050;
   wire FE_PHN4539_n1057;
   wire FE_PHN4538_n1034;
   wire FE_PHN4537_n2094;
   wire FE_PHN4536_n2307;
   wire FE_PHN4535_n1358;
   wire FE_PHN4534_n1229;
   wire FE_PHN4533_n1151;
   wire FE_PHN4532_n1552;
   wire FE_PHN4531_n1650;
   wire FE_PHN4530_n2388;
   wire FE_PHN4529_n1462;
   wire FE_PHN4528_n1135;
   wire FE_PHN4527_n1562;
   wire FE_PHN4526_n2191;
   wire FE_PHN4525_n943;
   wire FE_PHN4524_n1826;
   wire FE_PHN4523_n1035;
   wire FE_PHN4522_n1049;
   wire FE_PHN4521_n1386;
   wire FE_PHN4520_n1101;
   wire FE_PHN4519_n1345;
   wire FE_PHN4518_n1985;
   wire FE_PHN4517_n1879;
   wire FE_PHN4516_n1624;
   wire FE_PHN4515_n1379;
   wire FE_PHN4514_n1493;
   wire FE_PHN4513_n1728;
   wire FE_PHN4512_n1170;
   wire FE_PHN4511_n1468;
   wire FE_PHN4510_n1341;
   wire FE_PHN4509_n1201;
   wire FE_PHN4508_n1163;
   wire FE_PHN4507_n1169;
   wire FE_PHN4506_n1153;
   wire FE_PHN4505_n1936;
   wire FE_PHN4504_n1652;
   wire FE_PHN4503_n1278;
   wire FE_PHN4502_n1755;
   wire FE_PHN4501_n1084;
   wire FE_PHN4500_n1197;
   wire FE_PHN4499_n1008;
   wire FE_PHN4498_n1731;
   wire FE_PHN4497_n1950;
   wire FE_PHN4496_n912;
   wire FE_PHN4495_n1046;
   wire FE_PHN4494_n914;
   wire FE_PHN4493_n1376;
   wire FE_PHN4492_n1572;
   wire FE_PHN4491_n1974;
   wire FE_PHN4490_n1925;
   wire FE_PHN4489_n2311;
   wire FE_PHN4488_n1910;
   wire FE_PHN4487_n2159;
   wire FE_PHN4486_n1536;
   wire FE_PHN4485_n1234;
   wire FE_PHN4484_n1061;
   wire FE_PHN4483_n928;
   wire FE_PHN4482_n1325;
   wire FE_PHN4481_n927;
   wire FE_PHN4480_n1988;
   wire FE_PHN4479_n2238;
   wire FE_PHN4478_n1688;
   wire FE_PHN4477_n2301;
   wire FE_PHN4476_n1779;
   wire FE_PHN4475_n1865;
   wire FE_PHN4474_n1645;
   wire FE_PHN4473_n1312;
   wire FE_PHN4472_n1856;
   wire FE_PHN4471_n1089;
   wire FE_PHN4470_n1031;
   wire FE_PHN4469_n1592;
   wire FE_PHN4468_n1942;
   wire FE_PHN4467_n896;
   wire FE_PHN4466_n942;
   wire FE_PHN4465_n1014;
   wire FE_PHN4464_n1634;
   wire FE_PHN4463_n1628;
   wire FE_PHN4462_n2382;
   wire FE_PHN4461_n1514;
   wire FE_PHN4460_n1083;
   wire FE_PHN4459_n1993;
   wire FE_PHN4458_n2138;
   wire FE_PHN4457_n2322;
   wire FE_PHN4456_n1384;
   wire FE_PHN4455_n1588;
   wire FE_PHN4454_n1270;
   wire FE_PHN4453_n1122;
   wire FE_PHN4452_n2228;
   wire FE_PHN4451_n1683;
   wire FE_PHN4450_n2167;
   wire FE_PHN4449_n2149;
   wire FE_PHN4448_n2325;
   wire FE_PHN4447_n1047;
   wire FE_PHN4446_n1595;
   wire FE_PHN4445_n1635;
   wire FE_PHN4444_n1927;
   wire FE_PHN4443_n1568;
   wire FE_PHN4442_n2148;
   wire FE_PHN4441_n1269;
   wire FE_PHN4440_n1832;
   wire FE_PHN4439_n1076;
   wire FE_PHN4438_n1260;
   wire FE_PHN4437_n1969;
   wire FE_PHN4436_n1625;
   wire FE_PHN4435_n2232;
   wire FE_PHN4434_n1401;
   wire FE_PHN4433_n1373;
   wire FE_PHN4432_n1168;
   wire FE_PHN4431_n1295;
   wire FE_PHN4430_n945;
   wire FE_PHN4429_n1343;
   wire FE_PHN4428_n1432;
   wire FE_PHN4427_n1813;
   wire FE_PHN4426_n1540;
   wire FE_PHN4425_n1242;
   wire FE_PHN4424_n1166;
   wire FE_PHN4423_n1378;
   wire FE_PHN4422_n1971;
   wire FE_PHN4421_n2009;
   wire FE_PHN4420_n1853;
   wire FE_PHN4419_n1734;
   wire FE_PHN4418_n1056;
   wire FE_PHN4417_n2378;
   wire FE_PHN4416_n1286;
   wire FE_PHN4415_n1374;
   wire FE_PHN4414_n1094;
   wire FE_PHN4413_n1064;
   wire FE_PHN4412_n2306;
   wire FE_PHN4411_n1960;
   wire FE_PHN4410_n1955;
   wire FE_PHN4409_n956;
   wire FE_PHN4408_n2234;
   wire FE_PHN4407_n1573;
   wire FE_PHN4406_n1838;
   wire FE_PHN4405_n1298;
   wire FE_PHN4404_n921;
   wire FE_PHN4403_n1051;
   wire FE_PHN4402_n1603;
   wire FE_PHN4401_n1218;
   wire FE_PHN4400_n1140;
   wire FE_PHN4399_n1554;
   wire FE_PHN4398_n1368;
   wire FE_PHN4397_n2321;
   wire FE_PHN4396_n2387;
   wire FE_PHN4395_n983;
   wire FE_PHN4394_n1535;
   wire FE_PHN4393_n2267;
   wire FE_PHN4392_n1917;
   wire FE_PHN4391_n1265;
   wire FE_PHN4390_n1292;
   wire FE_PHN4389_n1478;
   wire FE_PHN4388_n1956;
   wire FE_PHN4387_n1530;
   wire FE_PHN4386_n1749;
   wire FE_PHN4385_n1892;
   wire FE_PHN4384_n2194;
   wire FE_PHN4383_n1288;
   wire FE_PHN4382_n963;
   wire FE_PHN4381_n1184;
   wire FE_PHN4380_n1464;
   wire FE_PHN4379_n1758;
   wire FE_PHN4378_n1776;
   wire FE_PHN4377_n1644;
   wire FE_PHN4376_n1767;
   wire FE_PHN4375_n2018;
   wire FE_PHN4374_n1160;
   wire FE_PHN4373_n1289;
   wire FE_PHN4372_n1217;
   wire FE_PHN4371_n1287;
   wire FE_PHN4370_n998;
   wire FE_PHN4369_n1240;
   wire FE_PHN4368_n1077;
   wire FE_PHN4367_n1097;
   wire FE_PHN4366_n1028;
   wire FE_PHN4365_n1953;
   wire FE_PHN4364_n1391;
   wire FE_PHN4363_n1351;
   wire FE_PHN4362_n1227;
   wire FE_PHN4361_n1377;
   wire FE_PHN4360_n1810;
   wire FE_PHN4359_n2174;
   wire FE_PHN4358_n2157;
   wire FE_PHN4357_n1016;
   wire FE_PHN4356_n1306;
   wire FE_PHN4355_n1675;
   wire FE_PHN4354_n1908;
   wire FE_PHN4353_n1697;
   wire FE_PHN4352_n1296;
   wire FE_PHN4351_n1366;
   wire FE_PHN4350_n1105;
   wire FE_PHN4349_n1560;
   wire FE_PHN4348_n2020;
   wire FE_PHN4347_n1861;
   wire FE_PHN4346_n2008;
   wire FE_PHN4345_n1964;
   wire FE_PHN4344_n1479;
   wire FE_PHN4343_n1342;
   wire FE_PHN4342_n1695;
   wire FE_PHN4341_n1275;
   wire FE_PHN4340_n1414;
   wire FE_PHN4339_n1946;
   wire FE_PHN4338_n1938;
   wire FE_PHN4337_n1238;
   wire FE_PHN4336_n975;
   wire FE_PHN4335_n1843;
   wire FE_PHN4334_n1461;
   wire FE_PHN4333_n2317;
   wire FE_PHN4332_n1670;
   wire FE_PHN4331_n2253;
   wire FE_PHN4330_n1791;
   wire FE_PHN4329_n2023;
   wire FE_PHN4328_n1060;
   wire FE_PHN4327_n1505;
   wire FE_PHN4326_n1633;
   wire FE_PHN4325_n929;
   wire FE_PHN4324_n1372;
   wire FE_PHN4323_n1859;
   wire FE_PHN4322_n2025;
   wire FE_PHN4321_n1301;
   wire FE_PHN4320_n1079;
   wire FE_PHN4319_n961;
   wire FE_PHN4318_n1396;
   wire FE_PHN4317_n1340;
   wire FE_PHN4316_n978;
   wire FE_PHN4315_n1305;
   wire FE_PHN4314_n1663;
   wire FE_PHN4313_n1648;
   wire FE_PHN4312_n1968;
   wire FE_PHN4311_n1096;
   wire FE_PHN4310_n1225;
   wire FE_PHN4309_n1346;
   wire FE_PHN4308_n1362;
   wire FE_PHN4307_n1104;
   wire FE_PHN4306_n1389;
   wire FE_PHN4305_n2013;
   wire FE_PHN4304_n2328;
   wire FE_PHN4303_n900;
   wire FE_PHN4302_n947;
   wire FE_PHN4301_n1222;
   wire FE_PHN4300_n1477;
   wire FE_PHN4299_n2029;
   wire FE_PHN4298_n2172;
   wire FE_PHN4297_n2258;
   wire FE_PHN4296_n1074;
   wire FE_PHN4295_n1082;
   wire FE_PHN4294_n976;
   wire FE_PHN4293_n1790;
   wire FE_PHN4292_n2027;
   wire FE_PHN4291_n1591;
   wire FE_PHN4290_n1845;
   wire FE_PHN4289_n1926;
   wire FE_PHN4288_n1700;
   wire FE_PHN4287_n1042;
   wire FE_PHN4286_n1280;
   wire FE_PHN4285_n2380;
   wire FE_PHN4284_n2065;
   wire FE_PHN4283_n1654;
   wire FE_PHN4282_n1816;
   wire FE_PHN4281_n1291;
   wire FE_PHN4280_n2239;
   wire FE_PHN4279_n2156;
   wire FE_PHN4278_n1963;
   wire FE_PHN4277_n916;
   wire FE_PHN4276_n1277;
   wire FE_PHN4275_n1279;
   wire FE_PHN4274_n2271;
   wire FE_PHN4273_n2111;
   wire FE_PHN4272_n2026;
   wire FE_PHN4271_n1931;
   wire FE_PHN4270_n1930;
   wire FE_PHN4269_n2323;
   wire FE_PHN4268_n1567;
   wire FE_PHN4267_n2115;
   wire FE_PHN4266_n2226;
   wire FE_PHN4265_n1496;
   wire FE_PHN4264_n1983;
   wire FE_PHN4263_n2329;
   wire FE_PHN4262_n1107;
   wire FE_PHN4261_n1991;
   wire FE_PHN4260_n2179;
   wire FE_PHN4259_n2140;
   wire FE_PHN4258_n2032;
   wire FE_PHN4257_n2207;
   wire FE_PHN4256_n934;
   wire FE_PHN4255_n1911;
   wire FE_PHN4254_n2184;
   wire FE_PHN4253_n1102;
   wire FE_PHN4252_n1081;
   wire FE_PHN4251_n1484;
   wire FE_PHN4250_n1881;
   wire FE_PHN4249_n1748;
   wire FE_PHN4248_n2012;
   wire FE_PHN4247_n1370;
   wire FE_PHN4246_n1017;
   wire FE_PHN4245_n1954;
   wire FE_PHN4244_n1445;
   wire FE_PHN4243_n1909;
   wire FE_PHN4242_n2280;
   wire FE_PHN4241_n1347;
   wire FE_PHN4240_n1236;
   wire FE_PHN4239_n1112;
   wire FE_PHN4238_n1784;
   wire FE_PHN4237_n1839;
   wire FE_PHN4236_n2045;
   wire FE_PHN4235_n1825;
   wire FE_PHN4234_n1054;
   wire FE_PHN4233_n952;
   wire FE_PHN4232_n1480;
   wire FE_PHN4231_n1574;
   wire FE_PHN4230_n1783;
   wire FE_PHN4229_n959;
   wire FE_PHN4228_n1765;
   wire FE_PHN4227_n1961;
   wire FE_PHN4226_n1040;
   wire FE_PHN4225_n1609;
   wire FE_PHN4224_n1707;
   wire FE_PHN4223_n1735;
   wire FE_PHN4222_n913;
   wire FE_PHN4221_n1780;
   wire FE_PHN4220_n2061;
   wire FE_PHN4219_n1590;
   wire FE_PHN4218_n1830;
   wire FE_PHN4217_n1257;
   wire FE_PHN4216_n1111;
   wire FE_PHN4215_n2189;
   wire FE_PHN4214_n1516;
   wire FE_PHN4213_n919;
   wire FE_PHN4212_n911;
   wire FE_PHN4211_n1510;
   wire FE_PHN4210_n1996;
   wire FE_PHN4209_n2123;
   wire FE_PHN4208_n1385;
   wire FE_PHN4207_n1995;
   wire FE_PHN4206_n2047;
   wire FE_PHN4205_n1841;
   wire FE_PHN4204_n1024;
   wire FE_PHN4203_n2151;
   wire FE_PHN4202_n2071;
   wire FE_PHN4201_n1751;
   wire FE_PHN4200_n1620;
   wire FE_PHN4199_n1837;
   wire FE_PHN4198_n1766;
   wire FE_PHN4197_n1668;
   wire FE_PHN4196_n2144;
   wire FE_PHN4195_n2318;
   wire FE_PHN4194_n1520;
   wire FE_PHN4193_n2052;
   wire FE_PHN4192_n970;
   wire FE_PHN4191_n1032;
   wire FE_PHN4190_n1885;
   wire FE_PHN4189_n2367;
   wire FE_PHN4188_n1828;
   wire FE_PHN4187_n1063;
   wire FE_PHN4186_n1418;
   wire FE_PHN4185_n1311;
   wire FE_PHN4184_n2287;
   wire FE_PHN4183_n1541;
   wire FE_PHN4182_n1407;
   wire FE_PHN4181_n1375;
   wire FE_PHN4180_n2038;
   wire FE_PHN4179_n2278;
   wire FE_PHN4178_n1504;
   wire FE_PHN4177_n1831;
   wire FE_PHN4176_n1250;
   wire FE_PHN4175_n1430;
   wire FE_PHN4174_n1455;
   wire FE_PHN4173_n1676;
   wire FE_PHN4172_n2040;
   wire FE_PHN4171_n1507;
   wire FE_PHN4170_n1161;
   wire FE_PHN4169_n2093;
   wire FE_PHN4168_n1958;
   wire FE_PHN4167_n1808;
   wire FE_PHN4166_n2163;
   wire FE_PHN4165_n1309;
   wire FE_PHN4164_n1124;
   wire FE_PHN4163_n2043;
   wire FE_PHN4162_n1742;
   wire FE_PHN4161_n1409;
   wire FE_PHN4160_n1420;
   wire FE_PHN4159_n1427;
   wire FE_PHN4158_n2222;
   wire FE_PHN4157_n1500;
   wire FE_PHN4156_n2241;
   wire FE_PHN4155_n2064;
   wire FE_PHN4154_n1937;
   wire FE_PHN4153_n1565;
   wire FE_PHN4152_n1545;
   wire FE_PHN4151_n1335;
   wire FE_PHN4150_n1330;
   wire FE_PHN4149_n1011;
   wire FE_PHN4148_n1677;
   wire FE_PHN4147_n979;
   wire FE_PHN4146_n933;
   wire FE_PHN4145_n1299;
   wire FE_PHN4144_n1900;
   wire FE_PHN4143_n1799;
   wire FE_PHN4142_n1449;
   wire FE_PHN4141_n1410;
   wire FE_PHN4140_n2147;
   wire FE_PHN4139_n971;
   wire FE_PHN4138_n1903;
   wire FE_PHN4137_n1320;
   wire FE_PHN4136_n1071;
   wire FE_PHN4135_n2289;
   wire FE_PHN4134_n984;
   wire FE_PHN4133_n2216;
   wire FE_PHN4132_n1665;
   wire FE_PHN4131_n1907;
   wire FE_PHN4130_n2131;
   wire FE_PHN4129_n1088;
   wire FE_PHN4128_n888;
   wire FE_PHN4127_n940;
   wire FE_PHN4126_n904;
   wire FE_PHN4125_n937;
   wire FE_PHN4124_n895;
   wire FE_PHN4123_n1773;
   wire FE_PHN4122_n1518;
   wire FE_PHN4121_n1851;
   wire FE_PHN4120_n2153;
   wire FE_PHN4119_n1716;
   wire FE_PHN4118_n2377;
   wire FE_PHN4117_n2303;
   wire FE_PHN4116_n1127;
   wire FE_PHN4115_n1254;
   wire FE_PHN4114_n1775;
   wire FE_PHN4113_n1469;
   wire FE_PHN4112_n1457;
   wire FE_PHN4111_n1923;
   wire FE_PHN4110_n1884;
   wire FE_PHN4109_n1777;
   wire FE_PHN4108_n1353;
   wire FE_PHN4107_n1782;
   wire FE_PHN4106_n2164;
   wire FE_PHN4105_n1788;
   wire FE_PHN4104_n1485;
   wire FE_PHN4103_n1337;
   wire FE_PHN4102_n1095;
   wire FE_PHN4101_n2248;
   wire FE_PHN4100_n1616;
   wire FE_PHN4099_n2128;
   wire FE_PHN4098_n1627;
   wire FE_PHN4097_n2331;
   wire FE_PHN4096_n1273;
   wire FE_PHN4095_n2039;
   wire FE_PHN4094_n1435;
   wire FE_PHN4093_n1606;
   wire FE_PHN4092_n1951;
   wire FE_PHN4091_n2291;
   wire FE_PHN4090_n1318;
   wire FE_PHN4089_n1513;
   wire FE_PHN4088_n2021;
   wire FE_PHN4087_n1333;
   wire FE_PHN4086_n1708;
   wire FE_PHN4085_n1471;
   wire FE_PHN4084_n1659;
   wire FE_PHN4083_n1920;
   wire FE_PHN4082_n1626;
   wire FE_PHN4081_n2236;
   wire FE_PHN4080_n1271;
   wire FE_PHN4079_n1336;
   wire FE_PHN4078_n2292;
   wire FE_PHN4077_n2240;
   wire FE_PHN4076_n1862;
   wire FE_PHN4075_n2003;
   wire FE_PHN4074_n968;
   wire FE_PHN4073_n1274;
   wire FE_PHN4072_n1196;
   wire FE_PHN4071_n1770;
   wire FE_PHN4070_n1792;
   wire FE_PHN4069_n1899;
   wire FE_PHN4068_n1334;
   wire FE_PHN4067_n2176;
   wire FE_PHN4066_n2002;
   wire FE_PHN4065_n1997;
   wire FE_PHN4064_n1736;
   wire FE_PHN4063_n2090;
   wire FE_PHN4062_n1975;
   wire FE_PHN4061_n1542;
   wire FE_PHN4060_n2221;
   wire FE_PHN4059_n1941;
   wire FE_PHN4058_n1395;
   wire FE_PHN4057_n991;
   wire FE_PHN4056_n1519;
   wire FE_PHN4055_n1725;
   wire FE_PHN4054_n2279;
   wire FE_PHN4053_n2000;
   wire FE_PHN4052_n1055;
   wire FE_PHN4051_n2122;
   wire FE_PHN4050_n2085;
   wire FE_PHN4049_n2063;
   wire FE_PHN4048_n890;
   wire FE_PHN4047_n1185;
   wire FE_PHN4046_n966;
   wire FE_PHN4045_n1578;
   wire FE_PHN4044_n1646;
   wire FE_PHN4043_n1740;
   wire FE_PHN4042_n1928;
   wire FE_PHN4041_n996;
   wire FE_PHN4040_n1023;
   wire FE_PHN4039_n950;
   wire FE_PHN4038_n1515;
   wire FE_PHN4037_n1466;
   wire FE_PHN4036_n1866;
   wire FE_PHN4035_n1544;
   wire FE_PHN4034_n2285;
   wire FE_PHN4033_n2101;
   wire FE_PHN4032_n1012;
   wire FE_PHN4031_n1403;
   wire FE_PHN4030_n1757;
   wire FE_PHN4029_n2100;
   wire FE_PHN4028_n2028;
   wire FE_PHN4027_n2386;
   wire FE_PHN4026_n1741;
   wire FE_PHN4025_n1128;
   wire FE_PHN4024_n986;
   wire FE_PHN4023_n1854;
   wire FE_PHN4022_n2281;
   wire FE_PHN4021_n2237;
   wire FE_PHN4020_n1547;
   wire FE_PHN4019_n1314;
   wire FE_PHN4018_n944;
   wire FE_PHN4017_n1456;
   wire FE_PHN4016_n1919;
   wire FE_PHN4015_n897;
   wire FE_PHN4014_n1297;
   wire FE_PHN4013_n1495;
   wire FE_PHN4012_n1600;
   wire FE_PHN4011_n2102;
   wire FE_PHN4010_n1143;
   wire FE_PHN4009_n2135;
   wire FE_PHN4008_n1474;
   wire FE_PHN4007_n1704;
   wire FE_PHN4006_n1522;
   wire FE_PHN4005_n2162;
   wire FE_PHN4004_n2048;
   wire FE_PHN4003_n894;
   wire FE_PHN4002_n1382;
   wire FE_PHN4001_n949;
   wire FE_PHN4000_n1875;
   wire FE_PHN3999_n1896;
   wire FE_PHN3998_n1890;
   wire FE_PHN3997_n2252;
   wire FE_PHN3996_n2096;
   wire FE_PHN3995_n2257;
   wire FE_PHN3994_n1310;
   wire FE_PHN3993_n1367;
   wire FE_PHN3992_n1175;
   wire FE_PHN3991_n2066;
   wire FE_PHN3990_n2268;
   wire FE_PHN3989_n1467;
   wire FE_PHN3988_n2262;
   wire FE_PHN3987_n1686;
   wire FE_PHN3986_n946;
   wire FE_PHN3985_n2127;
   wire FE_PHN3984_n1483;
   wire FE_PHN3983_n1844;
   wire FE_PHN3982_n2095;
   wire FE_PHN3981_n1850;
   wire FE_PHN3980_n1957;
   wire FE_PHN3979_n1948;
   wire FE_PHN3978_n972;
   wire FE_PHN3977_n903;
   wire FE_PHN3976_n982;
   wire FE_PHN3975_n1400;
   wire FE_PHN3974_n1846;
   wire FE_PHN3973_n1402;
   wire FE_PHN3972_n2110;
   wire FE_PHN3971_n1698;
   wire FE_PHN3970_n1680;
   wire FE_PHN3969_n1696;
   wire FE_PHN3968_n1664;
   wire FE_PHN3967_n1114;
   wire FE_PHN3966_n1433;
   wire FE_PHN3965_n1476;
   wire FE_PHN3964_n1715;
   wire FE_PHN3963_n905;
   wire FE_PHN3962_n1772;
   wire FE_PHN3961_n2006;
   wire FE_PHN3960_n1549;
   wire FE_PHN3959_n2108;
   wire FE_PHN3958_n2034;
   wire FE_PHN3957_n951;
   wire FE_PHN3956_n955;
   wire FE_PHN3955_n1709;
   wire FE_PHN3954_n2183;
   wire FE_PHN3953_n2211;
   wire FE_PHN3952_n1868;
   wire FE_PHN3951_n1913;
   wire FE_PHN3950_n1521;
   wire FE_PHN3949_n1576;
   wire FE_PHN3948_n1789;
   wire FE_PHN3947_n1316;
   wire FE_PHN3946_n1815;
   wire FE_PHN3945_n1821;
   wire FE_PHN3944_n2192;
   wire FE_PHN3943_n2272;
   wire FE_PHN3942_n922;
   wire FE_PHN3941_n985;
   wire FE_PHN3940_n1795;
   wire FE_PHN3939_n1000;
   wire FE_PHN3938_n1824;
   wire FE_PHN3937_n1747;
   wire FE_PHN3936_n2246;
   wire FE_PHN3935_n2109;
   wire FE_PHN3934_n1739;
   wire FE_PHN3933_n1580;
   wire FE_PHN3932_n1804;
   wire FE_PHN3931_n2249;
   wire FE_PHN3930_n2142;
   wire FE_PHN3929_n1802;
   wire FE_PHN3928_n1041;
   wire FE_PHN3927_n930;
   wire FE_PHN3926_n1869;
   wire FE_PHN3925_n1699;
   wire FE_PHN3924_n1524;
   wire FE_PHN3923_n2087;
   wire FE_PHN3922_n1397;
   wire FE_PHN3921_n1459;
   wire FE_PHN3920_n1441;
   wire FE_PHN3919_n967;
   wire FE_PHN3918_n1684;
   wire FE_PHN3917_n1921;
   wire FE_PHN3916_n2062;
   wire FE_PHN3915_n2168;
   wire FE_PHN3914_n2041;
   wire FE_PHN3913_n1858;
   wire FE_PHN3912_n1876;
   wire FE_PHN3911_n1428;
   wire FE_PHN3910_n1431;
   wire FE_PHN3909_n2001;
   wire FE_PHN3908_n2243;
   wire FE_PHN3907_n1491;
   wire FE_PHN3906_n1877;
   wire FE_PHN3905_n1883;
   wire FE_PHN3904_n1702;
   wire FE_PHN3903_n2143;
   wire FE_PHN3902_n1703;
   wire FE_PHN3901_n1711;
   wire FE_PHN3900_n2082;
   wire FE_PHN3899_n2118;
   wire FE_PHN3898_n2170;
   wire FE_PHN3897_n1448;
   wire FE_PHN3896_n1797;
   wire FE_PHN3895_n2051;
   wire FE_PHN3894_n1874;
   wire FE_PHN3893_n2286;
   wire FE_PHN3892_n1759;
   wire FE_PHN3891_n2072;
   wire FE_PHN3890_n1807;
   wire FE_PHN3889_n2077;
   wire FE_PHN3888_n2254;
   wire FE_PHN3887_n1701;
   wire FE_PHN3886_n2103;
   wire FE_PHN3885_n1768;
   wire FE_PHN3884_n923;
   wire FE_PHN3883_n1594;
   wire FE_PHN3882_n2230;
   wire FE_PHN3881_n1481;
   wire FE_PHN3880_n938;
   wire FE_PHN3879_n1497;
   wire FE_PHN3878_n1852;
   wire FE_PHN3877_n889;
   wire FE_PHN3876_n2205;
   wire FE_PHN3875_n1829;
   wire FE_PHN3874_n2244;
   wire FE_PHN3873_n2270;
   wire FE_PHN3872_n1778;
   wire FE_PHN3871_n1655;
   wire FE_PHN3870_n2208;
   wire FE_PHN3869_n962;
   wire FE_PHN3868_n1472;
   wire FE_PHN3867_n1762;
   wire FE_PHN3866_n908;
   wire FE_PHN3865_n1786;
   wire FE_PHN3864_n1738;
   wire FE_PHN3863_n2088;
   wire FE_PHN3862_n1743;
   wire FE_PHN3861_n2068;
   wire FE_PHN3860_n2173;
   wire FE_PHN3859_n1506;
   wire FE_PHN3858_n2374;
   wire FE_PHN3857_n1714;
   wire FE_PHN3856_n1998;
   wire FE_PHN3855_n1631;
   wire FE_PHN3854_n1710;
   wire FE_PHN3853_n964;
   wire FE_PHN3852_n2225;
   wire FE_PHN3851_n1691;
   wire FE_PHN3850_n1369;
   wire FE_PHN3849_n2245;
   wire FE_PHN3848_n2169;
   wire FE_PHN3847_n2199;
   wire FE_PHN3846_n1939;
   wire FE_PHN3845_n980;
   wire FE_PHN3844_n1498;
   wire FE_PHN3843_n2233;
   wire FE_PHN3842_n1499;
   wire FE_PHN3841_n1855;
   wire FE_PHN3840_n1523;
   wire FE_PHN3839_n1842;
   wire FE_PHN3838_n1417;
   wire FE_PHN3837_n1873;
   wire FE_PHN3836_n2132;
   wire FE_PHN3835_n1489;
   wire FE_PHN3834_n1490;
   wire FE_PHN3833_n1437;
   wire FE_PHN3832_n2075;
   wire FE_PHN3831_n2177;
   wire FE_PHN3830_n1593;
   wire FE_PHN3829_n1577;
   wire FE_PHN3828_n2203;
   wire FE_PHN3827_n1492;
   wire FE_PHN3826_n1870;
   wire FE_PHN3825_n1618;
   wire FE_PHN3824_n1835;
   wire FE_PHN3823_n2067;
   wire FE_PHN3822_n1894;
   wire FE_PHN3821_n1555;
   wire FE_PHN3820_n1415;
   wire FE_PHN3819_n2372;
   wire FE_PHN3818_n898;
   wire FE_PHN3817_n1745;
   wire FE_PHN3816_n1662;
   wire FE_PHN3815_n1880;
   wire FE_PHN3814_n2210;
   wire FE_PHN3813_n1672;
   wire FE_PHN3812_n1822;
   wire FE_PHN3811_n2265;
   wire FE_PHN3810_n1906;
   wire FE_PHN3809_n2269;
   wire FE_PHN3808_n1781;
   wire FE_PHN3807_n2214;
   wire FE_PHN3806_n2130;
   wire FE_PHN3805_n1673;
   wire FE_PHN3804_n2080;
   wire FE_PHN3803_n1473;
   wire FE_PHN3802_n2150;
   wire FE_PHN3801_n1502;
   wire FE_PHN3800_n1898;
   wire FE_PHN3799_n1723;
   wire FE_PHN3798_n1597;
   wire FE_PHN3797_n893;
   wire FE_PHN3796_n2086;
   wire FE_PHN3795_n1486;
   wire FE_PHN3794_n1604;
   wire FE_PHN3793_n1719;
   wire FE_PHN3792_n1438;
   wire FE_PHN3791_n2089;
   wire FE_PHN3790_n1817;
   wire FE_PHN3789_n1750;
   wire FE_PHN3788_n1399;
   wire FE_PHN3787_n1805;
   wire FE_PHN3786_n1945;
   wire FE_PHN3785_n2276;
   wire FE_PHN3784_n1657;
   wire FE_PHN3783_n2202;
   wire FE_PHN3782_n1364;
   wire FE_PHN3781_n1727;
   wire FE_PHN3780_n2213;
   wire FE_PHN3779_n1726;
   wire FE_PHN3778_n2079;
   wire FE_PHN3777_n2097;
   wire FE_PHN3776_n1660;
   wire FE_PHN3775_n1509;
   wire FE_PHN3774_n1967;
   wire FE_PHN3773_n1404;
   wire FE_PHN3772_n1756;
   wire FE_PHN3771_n1508;
   wire FE_PHN3770_n1860;
   wire FE_PHN3769_n1705;
   wire FE_PHN3768_n1729;
   wire FE_PHN3767_n1465;
   wire FE_PHN3766_n1882;
   wire FE_PHN3765_n2259;
   wire FE_PHN3764_n2083;
   wire FE_PHN3763_n2044;
   wire FE_PHN3762_n2055;
   wire FE_PHN3761_n1760;
   wire FE_PHN3760_n1671;
   wire FE_PHN3759_n1494;
   wire FE_PHN3758_n1871;
   wire FE_PHN3757_n1754;
   wire FE_PHN3756_n1443;
   wire FE_PHN3755_n1769;
   wire FE_PHN3754_n2198;
   wire FE_PHN3753_n1406;
   wire FE_PHN3752_n1798;
   wire FE_PHN3751_n2227;
   wire FE_PHN3750_n1801;
   wire FE_PHN3749_n1458;
   wire FE_PHN3748_n1787;
   wire FE_PHN3747_n1411;
   wire FE_PHN3746_n2178;
   wire FE_PHN3745_n2078;
   wire FE_PHN3744_n1803;
   wire FE_PHN3743_n2069;
   wire FE_PHN3742_n1451;
   wire FE_PHN3741_n2134;
   wire FE_PHN3740_n2242;
   wire FE_PHN3739_n2195;
   wire FE_PHN3738_n1863;
   wire FE_PHN3737_n2098;
   wire FE_PHN3736_n2264;
   wire FE_PHN3735_n1511;
   wire FE_PHN3734_n2054;
   wire FE_PHN3733_n1774;
   wire FE_PHN3732_n2260;
   wire FE_PHN3731_n1444;
   wire FE_PHN3730_n2187;
   wire FE_PHN3729_n2160;
   wire FE_PHN3728_n2251;
   wire FE_PHN3727_n2146;
   wire FE_PHN3726_n1823;
   wire FE_PHN3725_n2145;
   wire FE_PHN3724_n2218;
   wire FE_PHN3723_n1328;
   wire FE_PHN3722_n1840;
   wire FE_PHN3721_n1436;
   wire FE_PHN3720_n1752;
   wire FE_PHN3719_n1721;
   wire FE_PHN3718_n1429;
   wire FE_PHN3717_n2288;
   wire FE_PHN3716_n1439;
   wire FE_PHN3715_n2074;
   wire FE_PHN3714_n2217;
   wire FE_PHN3713_n1424;
   wire FE_PHN3712_n2112;
   wire FE_PHN3711_n2204;
   wire FE_PHN3710_n1656;
   wire FE_PHN3709_n1512;
   wire FE_PHN3708_n2099;
   wire FE_PHN3707_n2129;
   wire FE_PHN3706_n1694;
   wire FE_PHN3705_n2141;
   wire FE_PHN3704_n2224;
   wire FE_PHN3703_n2171;
   wire FE_PHN3702_n2106;
   wire FE_PHN3701_n2175;
   wire FE_PHN3700_n2107;
   wire FE_PHN3699_n1737;
   wire FE_PHN3698_n1722;
   wire FE_PHN3697_n1442;
   wire FE_PHN3696_n1849;
   wire FE_PHN3695_n2250;
   wire FE_PHN3694_n2196;
   wire FE_PHN3693_n2263;
   wire FE_PHN3692_n1667;
   wire FE_PHN3691_n2059;
   wire FE_PHN3690_n1864;
   wire FE_PHN3689_n1904;
   wire FE_PHN3688_n1487;
   wire FE_PHN3687_n1422;
   wire FE_PHN3686_n1814;
   wire FE_PHN3685_n1733;
   wire FE_PHN3684_n1463;
   wire FE_PHN3683_n1893;
   wire FE_PHN3682_n2200;
   wire FE_PHN3681_n1818;
   wire FE_PHN3680_n2206;
   wire FE_PHN3679_n1454;
   wire FE_PHN3678_n2057;
   wire FE_PHN3677_n2190;
   wire FE_PHN3676_n1692;
   wire FE_PHN3675_n1794;
   wire FE_PHN3674_n2092;
   wire FE_PHN3673_n2113;
   wire FE_PHN3672_n2136;
   wire FE_PHN3671_n1687;
   wire FE_PHN3670_n2050;
   wire FE_PHN3669_n1706;
   wire FE_PHN3668_n1452;
   wire FE_PHN3667_n1685;
   wire FE_PHN3666_n1446;
   wire FE_PHN3665_n1764;
   wire FE_PHN3664_n2070;
   wire FE_PHN3663_n2284;
   wire FE_PHN3662_n2158;
   wire FE_PHN3661_n1653;
   wire FE_PHN3660_n1503;
   wire FE_PHN3659_n1693;
   wire FE_PHN3658_n2056;
   wire FE_PHN3657_n2076;
   wire FE_PHN3656_n1833;
   wire FE_PHN3655_n2247;
   wire FE_PHN3654_n1834;
   wire FE_PHN3653_n2042;
   wire FE_PHN3652_n1679;
   wire FE_PHN3651_n1425;
   wire FE_PHN3650_n1412;
   wire FE_PHN3649_n1682;
   wire FE_PHN3648_n1678;
   wire FE_PHN3647_n1423;
   wire FE_PHN3646_n1994;
   wire FE_PHN3645_n1666;
   wire FE_PHN3644_n2152;
   wire FE_PHN3643_n1713;
   wire FE_PHN3642_n2105;
   wire FE_PHN3641_n1712;
   wire FE_PHN3640_n2073;
   wire FE_PHN3639_n2124;
   wire FE_PHN3638_n1405;
   wire FE_PHN3637_n2154;
   wire FE_PHN3636_n2220;
   wire FE_PHN3635_n2126;
   wire FE_PHN3634_n1848;
   wire FE_PHN3633_n1416;
   wire FE_PHN3632_n2231;
   wire FE_PHN3631_n1771;
   wire FE_PHN3630_n1720;
   wire FE_PHN3629_n2212;
   wire FE_PHN3628_n2193;
   wire FE_PHN3627_n2255;
   wire FE_PHN3626_n2235;
   wire FE_PHN3625_n1482;
   wire FE_PHN3624_n2266;
   wire FE_PHN3623_n1718;
   wire FE_PHN3622_n1450;
   wire FE_PHN3621_n2121;
   wire FE_PHN3620_n1658;
   wire FE_PHN3619_n1724;
   wire FE_PHN3618_n2215;
   wire FE_PHN3617_n2137;
   wire FE_PHN3616_n1717;
   wire FE_PHN3615_n1878;
   wire FE_PHN3614_n1891;
   wire FE_PHN3613_n1796;
   wire FE_PHN3612_n1763;
   wire FE_PHN3611_n1661;
   wire FE_PHN3444_key_mem_1407_;
   wire FE_PHN3437_key_mem_514_;
   wire FE_PHN3435_key_mem_1299_;
   wire FE_PHN3434_key_mem_898_;
   wire FE_PHN3433_key_mem_969_;
   wire FE_PHN3431_key_mem_1007_;
   wire FE_PHN3430_key_mem_394_;
   wire FE_PHN3429_key_mem_130_;
   wire FE_PHN3428_key_mem_138_;
   wire FE_PHN3427_key_mem_239_;
   wire FE_PHN3426_key_mem_1002_;
   wire FE_PHN3425_key_mem_409_;
   wire FE_PHN3424_key_mem_201_;
   wire FE_PHN3423_key_mem_234_;
   wire FE_PHN3422_key_mem_490_;
   wire FE_PHN3421_key_mem_874_;
   wire FE_PHN3420_key_mem_143_;
   wire FE_PHN3419_key_mem_1391_;
   wire FE_PHN3418_key_mem_255_;
   wire FE_PHN3417_key_mem_777_;
   wire FE_PHN3416_key_mem_522_;
   wire FE_PHN3415_key_mem_618_;
   wire FE_PHN3414_key_mem_585_;
   wire FE_PHN3413_key_mem_623_;
   wire FE_PHN3412_key_mem_770_;
   wire FE_PHN3411_key_mem_159_;
   wire FE_PHN3410_key_mem_543_;
   wire FE_PHN3409_n2430;
   wire FE_PHN3407_n883;
   wire FE_PHN3406_n881;
   wire FE_PHN3403_n2427;
   wire FE_PHN3373_n2868;
   wire FE_PHN3319_key_mem_1183_;
   wire FE_PHN3307_key_mem_1130_;
   wire FE_PHN3303_key_mem_1034_;
   wire FE_PHN3285_key_mem_1290_;
   wire FE_PHN3283_key_mem_15_;
   wire FE_PHN3275_key_mem_895_;
   wire FE_PHN3270_key_mem_889_;
   wire FE_PHN3258_key_mem_1393_;
   wire FE_PHN3248_key_mem_2_;
   wire FE_PHN3239_key_mem_1026_;
   wire FE_PHN3236_key_mem_879_;
   wire FE_PHN3234_key_mem_783_;
   wire FE_PHN3229_key_mem_1400_;
   wire FE_PHN3226_key_mem_386_;
   wire FE_PHN3221_key_mem_511_;
   wire FE_PHN3218_key_mem_403_;
   wire FE_PHN3215_key_mem_746_;
   wire FE_PHN3214_key_mem_665_;
   wire FE_PHN3213_key_mem_495_;
   wire FE_PHN3210_key_mem_799_;
   wire FE_PHN3209_key_mem_407_;
   wire FE_PHN3208_key_mem_127_;
   wire FE_PHN3207_key_mem_856_;
   wire FE_PHN3206_key_mem_10_;
   wire FE_PHN3205_key_mem_1289_;
   wire FE_PHN3204_key_mem_399_;
   wire FE_PHN3203_key_mem_863_;
   wire FE_PHN3201_key_mem_95_;
   wire FE_PHN3198_key_mem_791_;
   wire FE_PHN3197_key_mem_457_;
   wire FE_PHN3196_key_mem_761_;
   wire FE_PHN3195_key_mem_402_;
   wire FE_PHN3194_key_mem_18_;
   wire FE_PHN3189_key_mem_73_;
   wire FE_PHN3188_key_mem_19_;
   wire FE_PHN3187_key_mem_111_;
   wire FE_PHN3186_key_mem_841_;
   wire FE_PHN3185_key_mem_106_;
   wire FE_PHN3184_key_mem_415_;
   wire FE_PHN3094_key_mem_1303_;
   wire FE_PHN3091_key_mem_1279_;
   wire FE_PHN3089_key_mem_126_;
   wire FE_PHN3085_key_mem_31_;
   wire FE_PHN2855_n2423;
   wire FE_PHN2842_key_mem_1263_;
   wire FE_PHN2841_key_mem_1353_;
   wire FE_PHN2840_key_mem_1295_;
   wire FE_PHN2839_key_mem_1171_;
   wire FE_PHN2838_key_mem_1033_;
   wire FE_PHN2837_key_mem_1297_;
   wire FE_PHN2836_key_mem_1382_;
   wire FE_PHN2835_key_mem_1302_;
   wire FE_PHN2834_key_mem_1401_;
   wire FE_PHN2833_key_mem_1375_;
   wire FE_PHN2832_key_mem_650_;
   wire FE_PHN2831_key_mem_1262_;
   wire FE_PHN2830_key_mem_1368_;
   wire FE_PHN2829_key_mem_1305_;
   wire FE_PHN2828_key_mem_1351_;
   wire FE_PHN2827_key_mem_1304_;
   wire FE_PHN2826_key_mem_504_;
   wire FE_PHN2825_key_mem_1282_;
   wire FE_PHN2824_key_mem_753_;
   wire FE_PHN2823_key_mem_1298_;
   wire FE_PHN2820_n2421;
   wire FE_PHN2814_n880;
   wire FE_PHN2811_n2422;
   wire FE_PHN2810_key_mem_1386_;
   wire FE_PHN2799_n2391;
   wire FE_PHN2798_n2392;
   wire FE_PHN2795_n2390;
   wire FE_PHN2793_n2396;
   wire FE_PHN2792_n2395;
   wire FE_PHN2791_n2389;
   wire FE_PHN2790_n957;
   wire FE_PHN2789_key_mem_846_;
   wire FE_PHN2788_n918;
   wire FE_PHN2787_n1230;
   wire FE_PHN2786_n992;
   wire FE_PHN2785_n1329;
   wire FE_PHN2784_n935;
   wire FE_PHN2783_n1348;
   wire FE_PHN2782_n1355;
   wire FE_PHN2781_n1393;
   wire FE_PHN2780_n1371;
   wire FE_PHN2779_n965;
   wire FE_PHN2778_n973;
   wire FE_PHN2777_n886;
   wire FE_PHN2776_n1344;
   wire FE_PHN2775_n1294;
   wire FE_PHN2774_n1357;
   wire FE_PHN2773_n1319;
   wire FE_PHN2772_n931;
   wire FE_PHN2771_n1390;
   wire FE_PHN2770_n974;
   wire FE_PHN2769_n1075;
   wire FE_PHN2768_n1338;
   wire FE_PHN2767_n958;
   wire FE_PHN2766_n1363;
   wire FE_PHN2765_n1332;
   wire FE_PHN2764_n1380;
   wire FE_PHN2763_n1361;
   wire FE_PHN2762_n1356;
   wire FE_PHN2761_n1008;
   wire FE_PHN2760_n1387;
   wire FE_PHN2759_n1009;
   wire FE_PHN2758_n997;
   wire FE_PHN2757_n954;
   wire FE_PHN2756_n2188;
   wire FE_PHN2755_n2091;
   wire FE_PHN2754_n926;
   wire FE_PHN2753_n2229;
   wire FE_PHN2752_n1327;
   wire FE_PHN2751_n1340;
   wire FE_PHN2750_n1879;
   wire FE_PHN2749_n1298;
   wire FE_PHN2748_n1284;
   wire FE_PHN2747_n1744;
   wire FE_PHN2746_n1856;
   wire FE_PHN2745_n1272;
   wire FE_PHN2744_n1359;
   wire FE_PHN2743_n1368;
   wire FE_PHN2742_n932;
   wire FE_PHN2741_n1350;
   wire FE_PHN2740_n942;
   wire FE_PHN2739_n1339;
   wire FE_PHN2738_n885;
   wire FE_PHN2737_n1276;
   wire FE_PHN2736_n1269;
   wire FE_PHN2735_n1351;
   wire FE_PHN2734_n1286;
   wire FE_PHN2733_n1352;
   wire FE_PHN2732_n1315;
   wire FE_PHN2731_n939;
   wire FE_PHN2730_n1005;
   wire FE_PHN2729_n1307;
   wire FE_PHN2728_n2149;
   wire FE_PHN2727_n1501;
   wire FE_PHN2726_n1349;
   wire FE_PHN2725_n1384;
   wire FE_PHN2724_n1301;
   wire FE_PHN2723_n925;
   wire FE_PHN2722_n963;
   wire FE_PHN2721_n960;
   wire FE_PHN2720_n977;
   wire FE_PHN2719_n1358;
   wire FE_PHN2718_n1303;
   wire FE_PHN2717_n1468;
   wire FE_PHN2716_n1812;
   wire FE_PHN2715_n1392;
   wire FE_PHN2714_n1378;
   wire FE_PHN2713_n928;
   wire FE_PHN2712_n1001;
   wire FE_PHN2711_n1853;
   wire FE_PHN2710_n1278;
   wire FE_PHN2709_n1275;
   wire FE_PHN2708_n1377;
   wire FE_PHN2707_n2114;
   wire FE_PHN2706_n1341;
   wire FE_PHN2705_n1839;
   wire FE_PHN2704_n1293;
   wire FE_PHN2703_n993;
   wire FE_PHN2702_n899;
   wire FE_PHN2701_n1886;
   wire FE_PHN2700_n887;
   wire FE_PHN2699_n1372;
   wire FE_PHN2698_n937;
   wire FE_PHN2697_n2180;
   wire FE_PHN2696_n1109;
   wire FE_PHN2695_n1790;
   wire FE_PHN2694_n1292;
   wire FE_PHN2693_n2046;
   wire FE_PHN2692_n995;
   wire FE_PHN2691_n1302;
   wire FE_PHN2690_n915;
   wire FE_PHN2689_n1867;
   wire FE_PHN2688_n1330;
   wire FE_PHN2687_n1007;
   wire FE_PHN2686_n1383;
   wire FE_PHN2685_n999;
   wire FE_PHN2684_n929;
   wire FE_PHN2683_n1375;
   wire FE_PHN2682_n1432;
   wire FE_PHN2681_n1311;
   wire FE_PHN2680_n1346;
   wire FE_PHN2679_n1872;
   wire FE_PHN2678_n1281;
   wire FE_PHN2677_n2116;
   wire FE_PHN2676_n1836;
   wire FE_PHN2675_n896;
   wire FE_PHN2674_n1002;
   wire FE_PHN2673_n1347;
   wire FE_PHN2672_n1374;
   wire FE_PHN2671_n1493;
   wire FE_PHN2670_n2228;
   wire FE_PHN2669_n1765;
   wire FE_PHN2668_n2045;
   wire FE_PHN2667_n2119;
   wire FE_PHN2666_n1337;
   wire FE_PHN2665_n986;
   wire FE_PHN2664_n1746;
   wire FE_PHN2663_n1270;
   wire FE_PHN2662_n919;
   wire FE_PHN2661_n1810;
   wire FE_PHN2660_n998;
   wire FE_PHN2659_n1430;
   wire FE_PHN2658_n2060;
   wire FE_PHN2657_n914;
   wire FE_PHN2656_n1322;
   wire FE_PHN2655_n2038;
   wire FE_PHN2654_n1408;
   wire FE_PHN2653_n1324;
   wire FE_PHN2652_n940;
   wire FE_PHN2651_n1388;
   wire FE_PHN2650_n1479;
   wire FE_PHN2649_n2111;
   wire FE_PHN2648_n1516;
   wire FE_PHN2647_n1312;
   wire FE_PHN2646_n1271;
   wire FE_PHN2645_n2189;
   wire FE_PHN2644_n1427;
   wire FE_PHN2643_n1304;
   wire FE_PHN2642_n1784;
   wire FE_PHN2641_n907;
   wire FE_PHN2640_n989;
   wire FE_PHN2639_n1289;
   wire FE_PHN2638_n1758;
   wire FE_PHN2637_n1775;
   wire FE_PHN2636_n2234;
   wire FE_PHN2635_n1749;
   wire FE_PHN2634_n894;
   wire FE_PHN2633_n956;
   wire FE_PHN2632_n1277;
   wire FE_PHN2631_n1333;
   wire FE_PHN2630_n903;
   wire FE_PHN2629_n927;
   wire FE_PHN2628_n2249;
   wire FE_PHN2627_n1464;
   wire FE_PHN2626_n2223;
   wire FE_PHN2625_n1522;
   wire FE_PHN2624_n1300;
   wire FE_PHN2623_n1370;
   wire FE_PHN2622_n1813;
   wire FE_PHN2621_n2290;
   wire FE_PHN2620_n1888;
   wire FE_PHN2619_n1325;
   wire FE_PHN2618_n1517;
   wire FE_PHN2617_n1843;
   wire FE_PHN2616_n916;
   wire FE_PHN2615_n1309;
   wire FE_PHN2614_n945;
   wire FE_PHN2613_n1382;
   wire FE_PHN2612_n1663;
   wire FE_PHN2611_n1445;
   wire FE_PHN2610_n1291;
   wire FE_PHN2609_n911;
   wire FE_PHN2608_n2182;
   wire FE_PHN2607_n1859;
   wire FE_PHN2606_n1403;
   wire FE_PHN2605_n959;
   wire FE_PHN2604_n2287;
   wire FE_PHN2603_n1477;
   wire FE_PHN2602_n983;
   wire FE_PHN2601_n1816;
   wire FE_PHN2600_n2065;
   wire FE_PHN2599_n961;
   wire FE_PHN2598_n2039;
   wire FE_PHN2597_n2241;
   wire FE_PHN2596_n1793;
   wire FE_PHN2595_n1313;
   wire FE_PHN2594_n1316;
   wire FE_PHN2593_n1321;
   wire FE_PHN2592_n1455;
   wire FE_PHN2591_n1518;
   wire FE_PHN2590_n936;
   wire FE_PHN2589_n930;
   wire FE_PHN2588_n1394;
   wire FE_PHN2587_n910;
   wire FE_PHN2586_n1273;
   wire FE_PHN2585_n2109;
   wire FE_PHN2584_n1285;
   wire FE_PHN2583_n1279;
   wire FE_PHN2582_n1730;
   wire FE_PHN2581_n900;
   wire FE_PHN2580_n1369;
   wire FE_PHN2579_n2271;
   wire FE_PHN2578_n1435;
   wire FE_PHN2577_n1428;
   wire FE_PHN2576_n2176;
   wire FE_PHN2575_n1716;
   wire FE_PHN2574_n1362;
   wire FE_PHN2573_n2289;
   wire FE_PHN2572_n1676;
   wire FE_PHN2571_n1449;
   wire FE_PHN2570_n984;
   wire FE_PHN2569_n1700;
   wire FE_PHN2568_n949;
   wire FE_PHN2567_n1287;
   wire FE_PHN2566_n2166;
   wire FE_PHN2565_n943;
   wire FE_PHN2564_n970;
   wire FE_PHN2563_n934;
   wire FE_PHN2562_n1515;
   wire FE_PHN2561_n2094;
   wire FE_PHN2560_n2117;
   wire FE_PHN2559_n1689;
   wire FE_PHN2558_n1471;
   wire FE_PHN2557_n1353;
   wire FE_PHN2556_n988;
   wire FE_PHN2555_n933;
   wire FE_PHN2554_n1400;
   wire FE_PHN2553_n2084;
   wire FE_PHN2552_n2291;
   wire FE_PHN2551_n909;
   wire FE_PHN2550_n1838;
   wire FE_PHN2549_n1402;
   wire FE_PHN2548_n1011;
   wire FE_PHN2547_n2066;
   wire FE_PHN2546_n1703;
   wire FE_PHN2545_n905;
   wire FE_PHN2544_n1500;
   wire FE_PHN2543_n1874;
   wire FE_PHN2542_n1431;
   wire FE_PHN2541_n1708;
   wire FE_PHN2540_n967;
   wire FE_PHN2539_n1297;
   wire FE_PHN2538_n1824;
   wire FE_PHN2537_n2040;
   wire FE_PHN2536_n1809;
   wire FE_PHN2535_n2239;
   wire FE_PHN2534_n2139;
   wire FE_PHN2533_n2148;
   wire FE_PHN2532_n1485;
   wire FE_PHN2531_n1460;
   wire FE_PHN2530_n979;
   wire FE_PHN2529_n1695;
   wire FE_PHN2528_n1010;
   wire FE_PHN2527_n1318;
   wire FE_PHN2526_n2049;
   wire FE_PHN2525_n1495;
   wire FE_PHN2524_n2254;
   wire FE_PHN2523_n1699;
   wire FE_PHN2522_n1900;
   wire FE_PHN2521_n2253;
   wire FE_PHN2520_n2191;
   wire FE_PHN2519_n2115;
   wire FE_PHN2518_n1310;
   wire FE_PHN2517_n941;
   wire FE_PHN2516_n1761;
   wire FE_PHN2515_n1740;
   wire FE_PHN2514_n1686;
   wire FE_PHN2513_n1903;
   wire FE_PHN2512_n922;
   wire FE_PHN2511_n1326;
   wire FE_PHN2510_n1274;
   wire FE_PHN2509_n976;
   wire FE_PHN2508_n2232;
   wire FE_PHN2507_n898;
   wire FE_PHN2506_n2123;
   wire FE_PHN2505_n1776;
   wire FE_PHN2504_n2174;
   wire FE_PHN2503_n897;
   wire FE_PHN2502_n2248;
   wire FE_PHN2501_n1731;
   wire FE_PHN2500_n2230;
   wire FE_PHN2499_n2277;
   wire FE_PHN2498_n1861;
   wire FE_PHN2497_n1367;
   wire FE_PHN2496_n1670;
   wire FE_PHN2495_n980;
   wire FE_PHN2494_n1841;
   wire FE_PHN2493_n893;
   wire FE_PHN2492_n1478;
   wire FE_PHN2491_n1875;
   wire FE_PHN2490_n1884;
   wire FE_PHN2489_n921;
   wire FE_PHN2488_n2258;
   wire FE_PHN2487_n904;
   wire FE_PHN2486_n1842;
   wire FE_PHN2485_n1414;
   wire FE_PHN2484_n1725;
   wire FE_PHN2483_n1845;
   wire FE_PHN2482_n2072;
   wire FE_PHN2481_n996;
   wire FE_PHN2480_n912;
   wire FE_PHN2479_n982;
   wire FE_PHN2478_n1524;
   wire FE_PHN2477_n2037;
   wire FE_PHN2476_n2208;
   wire FE_PHN2475_n951;
   wire FE_PHN2474_n1897;
   wire FE_PHN2473_n1747;
   wire FE_PHN2472_n2150;
   wire FE_PHN2471_n2209;
   wire FE_PHN2470_n2118;
   wire FE_PHN2469_n1314;
   wire FE_PHN2468_n952;
   wire FE_PHN2467_n1795;
   wire FE_PHN2466_n2262;
   wire FE_PHN2465_n924;
   wire FE_PHN2464_n1701;
   wire FE_PHN2463_n1404;
   wire FE_PHN2462_n1857;
   wire FE_PHN2461_n1882;
   wire FE_PHN2460_n1000;
   wire FE_PHN2459_n1006;
   wire FE_PHN2458_n1334;
   wire FE_PHN2457_n889;
   wire FE_PHN2456_n2173;
   wire FE_PHN2455_n2275;
   wire FE_PHN2454_n1680;
   wire FE_PHN2453_n2103;
   wire FE_PHN2452_n2162;
   wire FE_PHN2451_n1806;
   wire FE_PHN2450_n1772;
   wire FE_PHN2449_n2135;
   wire FE_PHN2448_n1698;
   wire FE_PHN2447_n1892;
   wire FE_PHN2446_n1401;
   wire FE_PHN2445_n1328;
   wire FE_PHN2444_n1433;
   wire FE_PHN2443_n2108;
   wire FE_PHN2442_n1681;
   wire FE_PHN2441_n1434;
   wire FE_PHN2440_n901;
   wire FE_PHN2439_n2207;
   wire FE_PHN2438_n1822;
   wire FE_PHN2437_n1723;
   wire FE_PHN2436_n1735;
   wire FE_PHN2435_n1797;
   wire FE_PHN2434_n969;
   wire FE_PHN2433_n966;
   wire FE_PHN2432_n1780;
   wire FE_PHN2431_n950;
   wire FE_PHN2430_n1673;
   wire FE_PHN2429_n1821;
   wire FE_PHN2428_n1858;
   wire FE_PHN2427_n2051;
   wire FE_PHN2426_n1697;
   wire FE_PHN2425_n1748;
   wire FE_PHN2424_n2159;
   wire FE_PHN2423_n1707;
   wire FE_PHN2422_n1702;
   wire FE_PHN2421_n1831;
   wire FE_PHN2420_n1683;
   wire FE_PHN2419_n1830;
   wire FE_PHN2418_n938;
   wire FE_PHN2417_n895;
   wire FE_PHN2416_n1519;
   wire FE_PHN2415_n2276;
   wire FE_PHN2414_n1869;
   wire FE_PHN2413_n1837;
   wire FE_PHN2412_n2236;
   wire FE_PHN2411_n906;
   wire FE_PHN2410_n2043;
   wire FE_PHN2409_n1815;
   wire FE_PHN2408_n2184;
   wire FE_PHN2407_n1448;
   wire FE_PHN2406_n2161;
   wire FE_PHN2405_n964;
   wire FE_PHN2404_n1513;
   wire FE_PHN2403_n2087;
   wire FE_PHN2402_n1743;
   wire FE_PHN2401_n1398;
   wire FE_PHN2400_n1003;
   wire FE_PHN2399_n1484;
   wire FE_PHN2398_n1781;
   wire FE_PHN2397_n1783;
   wire FE_PHN2396_n1654;
   wire FE_PHN2395_n1483;
   wire FE_PHN2394_n1865;
   wire FE_PHN2393_n890;
   wire FE_PHN2392_n2153;
   wire FE_PHN2391_n1472;
   wire FE_PHN2390_n2134;
   wire FE_PHN2389_n1410;
   wire FE_PHN2388_n2216;
   wire FE_PHN2387_n2194;
   wire FE_PHN2386_n2269;
   wire FE_PHN2385_n1709;
   wire FE_PHN2384_n1474;
   wire FE_PHN2383_n1711;
   wire FE_PHN2382_n1870;
   wire FE_PHN2381_n2167;
   wire FE_PHN2380_n1458;
   wire FE_PHN2379_n2233;
   wire FE_PHN2378_n1466;
   wire FE_PHN2377_n2085;
   wire FE_PHN2376_n1502;
   wire FE_PHN2375_n1881;
   wire FE_PHN2374_n2226;
   wire FE_PHN2373_n1798;
   wire FE_PHN2372_n2075;
   wire FE_PHN2371_n1819;
   wire FE_PHN2370_n1694;
   wire FE_PHN2369_n1828;
   wire FE_PHN2368_n1899;
   wire FE_PHN2367_n2222;
   wire FE_PHN2366_n1755;
   wire FE_PHN2365_n1741;
   wire FE_PHN2364_n1421;
   wire FE_PHN2363_n2245;
   wire FE_PHN2362_n1465;
   wire FE_PHN2361_n2071;
   wire FE_PHN2360_n1742;
   wire FE_PHN2359_n2080;
   wire FE_PHN2358_n1523;
   wire FE_PHN2357_n2278;
   wire FE_PHN2356_n1504;
   wire FE_PHN2355_n2127;
   wire FE_PHN2354_n2130;
   wire FE_PHN2353_n1437;
   wire FE_PHN2352_n2227;
   wire FE_PHN2351_n2252;
   wire FE_PHN2350_n1674;
   wire FE_PHN2349_n1457;
   wire FE_PHN2348_n1719;
   wire FE_PHN2347_n2041;
   wire FE_PHN2346_n2270;
   wire FE_PHN2345_n2203;
   wire FE_PHN2344_n2113;
   wire FE_PHN2343_n1883;
   wire FE_PHN2342_n2128;
   wire FE_PHN2341_n2052;
   wire FE_PHN2340_n2102;
   wire FE_PHN2339_n2112;
   wire FE_PHN2338_n1893;
   wire FE_PHN2337_n1791;
   wire FE_PHN2336_n1794;
   wire FE_PHN2335_n1777;
   wire FE_PHN2334_n2156;
   wire FE_PHN2333_n2217;
   wire FE_PHN2332_n1811;
   wire FE_PHN2331_n1726;
   wire FE_PHN2330_n1778;
   wire FE_PHN2329_n2225;
   wire FE_PHN2328_n2213;
   wire FE_PHN2327_n1453;
   wire FE_PHN2326_n1514;
   wire FE_PHN2325_n2110;
   wire FE_PHN2324_n2053;
   wire FE_PHN2323_n1411;
   wire FE_PHN2322_n1512;
   wire FE_PHN2321_n1851;
   wire FE_PHN2320_n1901;
   wire FE_PHN2319_n2268;
   wire FE_PHN2318_n1767;
   wire FE_PHN2317_n1507;
   wire FE_PHN2316_n2244;
   wire FE_PHN2315_n1860;
   wire FE_PHN2314_n1684;
   wire FE_PHN2313_n1677;
   wire FE_PHN2312_n1475;
   wire FE_PHN2311_n1757;
   wire FE_PHN2310_n2177;
   wire FE_PHN2309_n1854;
   wire FE_PHN2308_n2086;
   wire FE_PHN2307_n2257;
   wire FE_PHN2306_n1728;
   wire FE_PHN2305_n1480;
   wire FE_PHN2304_n2292;
   wire FE_PHN2303_n1906;
   wire FE_PHN2302_n1436;
   wire FE_PHN2301_n2078;
   wire FE_PHN2300_n1469;
   wire FE_PHN2299_n1488;
   wire FE_PHN2298_n1409;
   wire FE_PHN2297_n1415;
   wire FE_PHN2296_n1441;
   wire FE_PHN2295_n1672;
   wire FE_PHN2294_n2074;
   wire FE_PHN2293_n2095;
   wire FE_PHN2292_n2238;
   wire FE_PHN2291_n1664;
   wire FE_PHN2290_n1454;
   wire FE_PHN2289_n1473;
   wire FE_PHN2288_n1399;
   wire FE_PHN2287_n2155;
   wire FE_PHN2286_n2272;
   wire FE_PHN2285_n1429;
   wire FE_PHN2284_n1876;
   wire FE_PHN2283_n2164;
   wire FE_PHN2282_n1770;
   wire FE_PHN2281_n1462;
   wire FE_PHN2280_n2101;
   wire FE_PHN2279_n2202;
   wire FE_PHN2278_n2145;
   wire FE_PHN2277_n1907;
   wire FE_PHN2276_n2093;
   wire FE_PHN2275_n2186;
   wire FE_PHN2274_n1508;
   wire FE_PHN2273_n1506;
   wire FE_PHN2272_n1467;
   wire FE_PHN2271_n1890;
   wire FE_PHN2270_n1682;
   wire FE_PHN2269_n2283;
   wire FE_PHN2268_n1662;
   wire FE_PHN2267_n1721;
   wire FE_PHN2266_n1823;
   wire FE_PHN2265_n1521;
   wire FE_PHN2264_n1503;
   wire FE_PHN2263_n1463;
   wire FE_PHN2262_n1443;
   wire FE_PHN2261_n2140;
   wire FE_PHN2260_n2201;
   wire FE_PHN2259_n1665;
   wire FE_PHN2258_n2240;
   wire FE_PHN2257_n2247;
   wire FE_PHN2256_n1801;
   wire FE_PHN2255_n1693;
   wire FE_PHN2254_n2100;
   wire FE_PHN2253_n2192;
   wire FE_PHN2252_n1756;
   wire FE_PHN2251_n2067;
   wire FE_PHN2250_n1862;
   wire FE_PHN2249_n1779;
   wire FE_PHN2248_n2131;
   wire FE_PHN2247_n2083;
   wire FE_PHN2246_n1685;
   wire FE_PHN2245_n2090;
   wire FE_PHN2244_n2097;
   wire FE_PHN2243_n1866;
   wire FE_PHN2242_n1817;
   wire FE_PHN2241_n2220;
   wire FE_PHN2240_n1792;
   wire FE_PHN2239_n2055;
   wire FE_PHN2238_n1720;
   wire FE_PHN2237_n1509;
   wire FE_PHN2236_n1787;
   wire FE_PHN2235_n1727;
   wire FE_PHN2234_n1889;
   wire FE_PHN2233_n1788;
   wire FE_PHN2232_n1785;
   wire FE_PHN2231_n2165;
   wire FE_PHN2230_n1868;
   wire FE_PHN2229_n1877;
   wire FE_PHN2228_n1451;
   wire FE_PHN2227_n2126;
   wire FE_PHN2226_n2224;
   wire FE_PHN2225_n2255;
   wire FE_PHN2224_n1456;
   wire FE_PHN2223_n1494;
   wire FE_PHN2222_n2274;
   wire FE_PHN2221_n1803;
   wire FE_PHN2220_n2219;
   wire FE_PHN2219_n1754;
   wire FE_PHN2218_n1898;
   wire FE_PHN2217_n2154;
   wire FE_PHN2216_n2250;
   wire FE_PHN2215_n2260;
   wire FE_PHN2214_n1863;
   wire FE_PHN2213_n1696;
   wire FE_PHN2212_n1844;
   wire FE_PHN2211_n2178;
   wire FE_PHN2210_n1832;
   wire FE_PHN2209_n2231;
   wire FE_PHN2208_n2195;
   wire FE_PHN2207_n1840;
   wire FE_PHN2206_n1444;
   wire FE_PHN2205_n1492;
   wire FE_PHN2204_n2129;
   wire FE_PHN2203_n1871;
   wire FE_PHN2202_n2082;
   wire FE_PHN2201_n2193;
   wire FE_PHN2200_n1440;
   wire FE_PHN2199_n2059;
   wire FE_PHN2198_n1679;
   wire FE_PHN2197_n1729;
   wire FE_PHN2196_n1834;
   wire FE_PHN2195_n2256;
   wire FE_PHN2194_n2285;
   wire FE_PHN2193_n2261;
   wire FE_PHN2192_n1804;
   wire FE_PHN2191_n1482;
   wire FE_PHN2190_n1420;
   wire FE_PHN2189_n1905;
   wire FE_PHN2188_n2054;
   wire FE_PHN2187_n2120;
   wire FE_PHN2186_n2197;
   wire FE_PHN2185_n1820;
   wire FE_PHN2184_n2242;
   wire FE_PHN2183_n1760;
   wire FE_PHN2182_n2282;
   wire FE_PHN2181_n1773;
   wire FE_PHN2180_n2136;
   wire FE_PHN2179_n1497;
   wire FE_PHN2178_n2212;
   wire FE_PHN2177_n2200;
   wire FE_PHN2176_n2288;
   wire FE_PHN2175_n1722;
   wire FE_PHN2174_n1847;
   wire FE_PHN2173_n1827;
   wire FE_PHN2172_n1705;
   wire FE_PHN2171_n1864;
   wire FE_PHN2170_n1446;
   wire FE_PHN2169_n1789;
   wire FE_PHN2168_n2190;
   wire FE_PHN2167_n1669;
   wire FE_PHN2166_n1759;
   wire FE_PHN2165_n1715;
   wire FE_PHN2164_n1406;
   wire FE_PHN2163_n1887;
   wire FE_PHN2162_n2070;
   wire FE_PHN2161_n2181;
   wire FE_PHN2160_n1850;
   wire FE_PHN2159_n2210;
   wire FE_PHN2158_n1904;
   wire FE_PHN2157_n2099;
   wire FE_PHN2156_n1714;
   wire FE_PHN2155_n2096;
   wire FE_PHN2154_n1489;
   wire FE_PHN2153_n1724;
   wire FE_PHN2152_n2163;
   wire FE_PHN2151_n1704;
   wire FE_PHN2150_n1774;
   wire FE_PHN2149_n1835;
   wire FE_PHN2148_n1848;
   wire FE_PHN2147_n2204;
   wire FE_PHN2146_n2237;
   wire FE_PHN2145_n2142;
   wire FE_PHN2144_n2160;
   wire FE_PHN2143_n1802;
   wire FE_PHN2142_n1656;
   wire FE_PHN2141_n1397;
   wire FE_PHN2140_n2175;
   wire FE_PHN2139_n2273;
   wire FE_PHN2138_n2121;
   wire FE_PHN2137_n2206;
   wire FE_PHN2136_n1825;
   wire FE_PHN2135_n1653;
   wire FE_PHN2134_n1846;
   wire FE_PHN2133_n1424;
   wire FE_PHN2132_n2141;
   wire FE_PHN2131_n1442;
   wire FE_PHN2130_n1849;
   wire FE_PHN2129_n2137;
   wire FE_PHN2128_n1733;
   wire FE_PHN2127_n2081;
   wire FE_PHN2126_n2196;
   wire FE_PHN2125_n1894;
   wire FE_PHN2124_n1452;
   wire FE_PHN2123_n2218;
   wire FE_PHN2122_n1718;
   wire FE_PHN2121_n1486;
   wire FE_PHN2120_n1692;
   wire FE_PHN2119_n2259;
   wire FE_PHN2118_n1878;
   wire FE_PHN2117_n1826;
   wire FE_PHN2116_n1690;
   wire FE_PHN2115_n2132;
   wire FE_PHN2114_n2251;
   wire FE_PHN2113_n2146;
   wire FE_PHN2112_n1491;
   wire FE_PHN2111_n1818;
   wire FE_PHN2110_n1880;
   wire FE_PHN2109_n2158;
   wire FE_PHN2108_n2068;
   wire FE_PHN2107_n1450;
   wire FE_PHN2106_n1666;
   wire FE_PHN2105_n1852;
   wire FE_PHN2104_n1417;
   wire FE_PHN2103_n1487;
   wire FE_PHN2102_n1713;
   wire FE_PHN2101_n2062;
   wire FE_PHN2100_n1717;
   wire FE_PHN2099_n1855;
   wire FE_PHN2098_n1422;
   wire FE_PHN2097_n1891;
   wire FE_PHN2096_n1814;
   wire FE_PHN2095_n1426;
   wire FE_PHN2094_n2168;
   wire FE_PHN2093_n2215;
   wire FE_PHN2092_n1833;
   wire FE_PHN2091_n1407;
   wire FE_PHN2090_n2152;
   wire FE_PHN2089_n1706;
   wire FE_PHN2088_n2284;
   wire FE_PHN2087_n1425;
   wire FE_PHN2086_n2198;
   wire FE_PHN2085_n1405;
   wire FE_PHN2084_n2079;
   wire FE_PHN2083_n2214;
   wire FE_PHN2082_n1412;
   wire FE_PHN2081_n1710;
   wire FE_PHN2080_n1499;
   wire FE_PHN2079_n1496;
   wire FE_PHN2078_n1873;
   wire FE_PHN2077_n1423;
   wire FE_PHN2076_n2105;
   wire FE_PHN2075_n1762;
   wire FE_PHN2074_n2089;
   wire FE_PHN2073_n1678;
   wire FE_PHN2072_n2286;
   wire FE_PHN2071_n2138;
   wire FE_PHN2070_n2211;
   wire FE_PHN2069_n1829;
   wire FE_PHN2068_n1753;
   wire FE_PHN2067_n2243;
   wire FE_PHN2066_n1498;
   wire FE_PHN2065_n1796;
   wire FE_PHN2064_n2246;
   wire FE_PHN2063_n1712;
   wire FE_PHN2062_n1661;
   wire FE_PHN2061_n1691;
   wire FE_PHN2060_n1490;
   wire FE_PHN2059_n1459;
   wire FE_PHN2058_n2199;
   wire FE_PHN2057_n2088;
   wire FE_PHN2056_n1764;
   wire FE_PHN2055_n1763;
   wire FE_PHN2054_n1771;
   wire FE_PHN2053_n2044;
   wire FE_PHN2052_n2221;
   wire FE_PHN2051_n1805;
   wire FE_PHN2050_n1687;
   wire FE_PHN2049_n1885;
   wire FE_PHN2048_n2235;
   wire FE_PHN2047_n2104;
   wire FE_PHN2046_n1416;
   wire FE_PHN2045_n2073;
   wire FE_PHN2044_n1732;
   wire FE_PHN2043_n1769;
   wire FE_PHN2042_n2069;
   wire FE_PHN2041_n2098;
   wire FE_PHN2040_n2092;
   wire FE_PHN2039_n1511;
   wire FE_PHN2038_n2393;
   wire FE_PHN2036_n2394;
   wire FE_PHN2009_n1799;
   wire FE_PHN2008_n1786;
   wire FE_PHN2007_keymem_sboxw_13_;
   wire FE_PHN2006_keymem_sboxw_5_;
   wire FE_PHN2005_keymem_sboxw_20_;
   wire FE_PHN2004_keymem_sboxw_12_;
   wire FE_PHN2003_keymem_sboxw_4_;
   wire FE_PHN2002_keymem_sboxw_11_;
   wire FE_PHN2001_keymem_sboxw_8_;
   wire FE_PHN2000_keymem_sboxw_3_;
   wire FE_PHN1998_keymem_sboxw_17_;
   wire FE_PHN1997_keymem_sboxw_16_;
   wire FE_PHN1992_keymem_sboxw_19_;
   wire FE_PHN1991_keymem_sboxw_9_;
   wire FE_PHN1989_rcon_reg_6_;
   wire FE_PHN1974_keymem_sboxw_14_;
   wire FE_PHN1972_keymem_sboxw_15_;
   wire FE_PHN1969_keymem_sboxw_23_;
   wire FE_PHN1965_keymem_sboxw_22_;
   wire FE_PHN1962_keymem_sboxw_10_;
   wire FE_PHN1959_keymem_sboxw_0_;
   wire FE_PHN1958_keymem_sboxw_18_;
   wire FE_PHN1957_keymem_sboxw_1_;
   wire FE_PHN1930_key_mem_1082_;
   wire FE_PHN1917_key_mem_1207_;
   wire FE_PHN1905_key_mem_1046_;
   wire FE_PHN1899_key_mem_1272_;
   wire FE_PHN1894_key_mem_1044_;
   wire FE_PHN1893_key_mem_1101_;
   wire FE_PHN1892_key_mem_1029_;
   wire FE_PHN1891_key_mem_1068_;
   wire FE_PHN1889_key_mem_1071_;
   wire FE_PHN1888_key_mem_1039_;
   wire FE_PHN1887_key_mem_1100_;
   wire FE_PHN1885_key_mem_1114_;
   wire FE_PHN1884_key_mem_1151_;
   wire FE_PHN1883_key_mem_1153_;
   wire FE_PHN1882_key_mem_1025_;
   wire FE_PHN1881_key_mem_1040_;
   wire FE_PHN1880_key_mem_1045_;
   wire FE_PHN1879_key_mem_688_;
   wire FE_PHN1878_n1167;
   wire FE_PHN1877_key_mem_1255_;
   wire FE_PHN1876_key_mem_1049_;
   wire FE_PHN1874_key_mem_1143_;
   wire FE_PHN1873_key_mem_1061_;
   wire FE_PHN1872_key_mem_1060_;
   wire FE_PHN1871_key_mem_1106_;
   wire FE_PHN1870_key_mem_1138_;
   wire FE_PHN1869_key_mem_1088_;
   wire FE_PHN1868_key_mem_1053_;
   wire FE_PHN1867_key_mem_1069_;
   wire FE_PHN1866_key_mem_1078_;
   wire FE_PHN1864_key_mem_1055_;
   wire FE_PHN1863_key_mem_1094_;
   wire FE_PHN1862_key_mem_1030_;
   wire FE_PHN1861_key_mem_1072_;
   wire FE_PHN1860_key_mem_1112_;
   wire FE_PHN1859_key_mem_1099_;
   wire FE_PHN1858_key_mem_1144_;
   wire FE_PHN1857_key_mem_1083_;
   wire FE_PHN1856_key_mem_1085_;
   wire FE_PHN1855_key_mem_1103_;
   wire FE_PHN1854_key_mem_1127_;
   wire FE_PHN1853_key_mem_1028_;
   wire FE_PHN1852_key_mem_1064_;
   wire FE_PHN1851_key_mem_349_;
   wire FE_PHN1850_key_mem_1121_;
   wire FE_PHN1849_key_mem_376_;
   wire FE_PHN1848_key_mem_647_;
   wire FE_PHN1847_n1162;
   wire FE_PHN1846_key_mem_1142_;
   wire FE_PHN1844_key_mem_352_;
   wire FE_PHN1843_key_mem_1116_;
   wire FE_PHN1841_key_mem_1092_;
   wire FE_PHN1840_key_mem_1041_;
   wire FE_PHN1839_key_mem_1059_;
   wire FE_PHN1837_n2267;
   wire FE_PHN1835_key_mem_1084_;
   wire FE_PHN1834_key_mem_1311_;
   wire FE_PHN1833_key_mem_1043_;
   wire FE_PHN1832_key_mem_1057_;
   wire FE_PHN1831_key_mem_724_;
   wire FE_PHN1830_key_mem_1090_;
   wire FE_PHN1829_key_mem_1079_;
   wire FE_PHN1828_key_mem_755_;
   wire FE_PHN1827_n1181;
   wire FE_PHN1826_key_mem_334_;
   wire FE_PHN1824_key_mem_738_;
   wire FE_PHN1823_key_mem_1115_;
   wire FE_PHN1822_key_mem_1133_;
   wire FE_PHN1821_key_mem_1104_;
   wire FE_PHN1820_key_mem_713_;
   wire FE_PHN1819_key_mem_1140_;
   wire FE_PHN1818_key_mem_1113_;
   wire FE_PHN1817_key_mem_1119_;
   wire FE_PHN1816_key_mem_1128_;
   wire FE_PHN1814_key_mem_1150_;
   wire FE_PHN1813_key_mem_1066_;
   wire FE_PHN1812_n1595;
   wire FE_PHN1811_key_mem_1036_;
   wire FE_PHN1810_key_mem_1136_;
   wire FE_PHN1809_key_mem_644_;
   wire FE_PHN1808_key_mem_1148_;
   wire FE_PHN1807_key_mem_360_;
   wire FE_PHN1806_key_mem_318_;
   wire FE_PHN1805_key_mem_1147_;
   wire FE_PHN1804_key_mem_737_;
   wire FE_PHN1803_key_mem_1118_;
   wire FE_PHN1802_key_mem_285_;
   wire FE_PHN1801_n1240;
   wire FE_PHN1800_key_mem_1191_;
   wire FE_PHN1799_key_mem_1097_;
   wire FE_PHN1798_key_mem_1076_;
   wire FE_PHN1797_key_mem_661_;
   wire FE_PHN1796_n1579;
   wire FE_PHN1795_key_mem_311_;
   wire FE_PHN1794_key_mem_709_;
   wire FE_PHN1793_key_mem_353_;
   wire FE_PHN1792_key_mem_1169_;
   wire FE_PHN1791_key_mem_1135_;
   wire FE_PHN1790_key_mem_1093_;
   wire FE_PHN1789_key_mem_1077_;
   wire FE_PHN1788_key_mem_1037_;
   wire FE_PHN1787_key_mem_1109_;
   wire FE_PHN1786_key_mem_1134_;
   wire FE_PHN1785_key_mem_302_;
   wire FE_PHN1784_key_mem_1051_;
   wire FE_PHN1783_key_mem_1081_;
   wire FE_PHN1782_n2179;
   wire FE_PHN1781_key_mem_1123_;
   wire FE_PHN1780_key_mem_1267_;
   wire FE_PHN1779_key_mem_694_;
   wire FE_PHN1778_key_mem_1095_;
   wire FE_PHN1777_key_mem_1132_;
   wire FE_PHN1776_key_mem_684_;
   wire FE_PHN1775_key_mem_344_;
   wire FE_PHN1774_n1266;
   wire FE_PHN1773_key_mem_1074_;
   wire FE_PHN1772_key_mem_1050_;
   wire FE_PHN1771_key_mem_696_;
   wire FE_PHN1770_key_mem_723_;
   wire FE_PHN1769_key_mem_1054_;
   wire FE_PHN1768_n2047;
   wire FE_PHN1767_n1257;
   wire FE_PHN1766_key_mem_1278_;
   wire FE_PHN1765_key_mem_764_;
   wire FE_PHN1764_key_mem_1137_;
   wire FE_PHN1763_key_mem_689_;
   wire FE_PHN1762_key_mem_1145_;
   wire FE_PHN1761_key_mem_1047_;
   wire FE_PHN1760_key_mem_1031_;
   wire FE_PHN1759_n1668;
   wire FE_PHN1758_key_mem_1070_;
   wire FE_PHN1757_key_mem_359_;
   wire FE_PHN1756_key_mem_1098_;
   wire FE_PHN1755_key_mem_708_;
   wire FE_PHN1754_key_mem_351_;
   wire FE_PHN1752_n1168;
   wire FE_PHN1751_key_mem_758_;
   wire FE_PHN1750_key_mem_707_;
   wire FE_PHN1749_key_mem_675_;
   wire FE_PHN1748_key_mem_1141_;
   wire FE_PHN1747_key_mem_682_;
   wire FE_PHN1746_key_mem_732_;
   wire FE_PHN1745_key_mem_1105_;
   wire FE_PHN1744_key_mem_659_;
   wire FE_PHN1743_key_mem_1058_;
   wire FE_PHN1742_key_mem_328_;
   wire FE_PHN1740_key_mem_1120_;
   wire FE_PHN1739_key_mem_345_;
   wire FE_PHN1738_key_mem_260_;
   wire FE_PHN1737_n1895;
   wire FE_PHN1736_n1596;
   wire FE_PHN1735_key_mem_291_;
   wire FE_PHN1734_key_mem_1152_;
   wire FE_PHN1733_n1547;
   wire FE_PHN1732_n1751;
   wire FE_PHN1731_key_mem_693_;
   wire FE_PHN1730_key_mem_1080_;
   wire FE_PHN1729_key_mem_297_;
   wire FE_PHN1728_n2185;
   wire FE_PHN1727_key_mem_269_;
   wire FE_PHN1726_key_mem_374_;
   wire FE_PHN1725_key_mem_348_;
   wire FE_PHN1724_key_mem_660_;
   wire FE_PHN1723_key_mem_759_;
   wire FE_PHN1722_key_mem_648_;
   wire FE_PHN1721_key_mem_704_;
   wire FE_PHN1720_key_mem_1188_;
   wire FE_PHN1719_key_mem_1042_;
   wire FE_PHN1718_key_mem_721_;
   wire FE_PHN1717_key_mem_309_;
   wire FE_PHN1716_key_mem_324_;
   wire FE_PHN1715_key_mem_279_;
   wire FE_PHN1714_key_mem_341_;
   wire FE_PHN1713_key_mem_1032_;
   wire FE_PHN1712_key_mem_1075_;
   wire FE_PHN1711_key_mem_256_;
   wire FE_PHN1710_key_mem_316_;
   wire FE_PHN1709_n1258;
   wire FE_PHN1708_n1734;
   wire FE_PHN1707_key_mem_343_;
   wire FE_PHN1706_key_mem_671_;
   wire FE_PHN1705_n2143;
   wire FE_PHN1703_key_mem_258_;
   wire FE_PHN1702_key_mem_710_;
   wire FE_PHN1701_key_mem_1089_;
   wire FE_PHN1700_key_mem_1215_;
   wire FE_PHN1699_key_mem_262_;
   wire FE_PHN1698_key_mem_698_;
   wire FE_PHN1697_key_mem_266_;
   wire FE_PHN1696_key_mem_680_;
   wire FE_PHN1695_key_mem_716_;
   wire FE_PHN1694_key_mem_673_;
   wire FE_PHN1693_n1578;
   wire FE_PHN1692_key_mem_739_;
   wire FE_PHN1691_key_mem_308_;
   wire FE_PHN1690_key_mem_346_;
   wire FE_PHN1689_key_mem_325_;
   wire FE_PHN1688_key_mem_265_;
   wire FE_PHN1687_key_mem_662_;
   wire FE_PHN1686_n1438;
   wire FE_PHN1685_n1896;
   wire FE_PHN1684_key_mem_288_;
   wire FE_PHN1683_key_mem_323_;
   wire FE_PHN1682_key_mem_263_;
   wire FE_PHN1681_n1552;
   wire FE_PHN1680_key_mem_734_;
   wire FE_PHN1679_key_mem_757_;
   wire FE_PHN1678_key_mem_715_;
   wire FE_PHN1677_key_mem_363_;
   wire FE_PHN1676_n1581;
   wire FE_PHN1675_n1655;
   wire FE_PHN1674_n2172;
   wire FE_PHN1673_n1807;
   wire FE_PHN1672_key_mem_272_;
   wire FE_PHN1671_key_mem_731_;
   wire FE_PHN1670_key_mem_380_;
   wire FE_PHN1669_n2077;
   wire FE_PHN1668_key_mem_742_;
   wire FE_PHN1667_key_mem_322_;
   wire FE_PHN1666_key_mem_730_;
   wire FE_PHN1665_n2205;
   wire FE_PHN1664_n1461;
   wire FE_PHN1663_key_mem_687_;
   wire FE_PHN1662_n1539;
   wire FE_PHN1661_key_mem_677_;
   wire FE_PHN1660_key_mem_663_;
   wire FE_PHN1659_key_mem_354_;
   wire FE_PHN1658_key_mem_317_;
   wire FE_PHN1657_key_mem_656_;
   wire FE_PHN1656_key_mem_701_;
   wire FE_PHN1655_key_mem_358_;
   wire FE_PHN1654_n1531;
   wire FE_PHN1653_key_mem_342_;
   wire FE_PHN1652_key_mem_261_;
   wire FE_PHN1651_n2169;
   wire FE_PHN1650_key_mem_301_;
   wire FE_PHN1649_n1671;
   wire FE_PHN1648_n2280;
   wire FE_PHN1647_n1520;
   wire FE_PHN1646_key_mem_726_;
   wire FE_PHN1645_key_mem_697_;
   wire FE_PHN1644_key_mem_370_;
   wire FE_PHN1643_n1675;
   wire FE_PHN1642_key_mem_728_;
   wire FE_PHN1641_key_mem_674_;
   wire FE_PHN1640_n1745;
   wire FE_PHN1639_key_mem_274_;
   wire FE_PHN1638_key_mem_692_;
   wire FE_PHN1637_key_mem_338_;
   wire FE_PHN1636_key_mem_750_;
   wire FE_PHN1635_key_mem_315_;
   wire FE_PHN1634_key_mem_280_;
   wire FE_PHN1633_key_mem_307_;
   wire FE_PHN1632_key_mem_264_;
   wire FE_PHN1631_key_mem_756_;
   wire FE_PHN1630_key_mem_685_;
   wire FE_PHN1629_n2151;
   wire FE_PHN1628_n2125;
   wire FE_PHN1627_key_mem_329_;
   wire FE_PHN1626_key_mem_270_;
   wire FE_PHN1625_n1618;
   wire FE_PHN1624_key_mem_645_;
   wire FE_PHN1623_key_mem_281_;
   wire FE_PHN1622_key_mem_278_;
   wire FE_PHN1621_key_mem_321_;
   wire FE_PHN1620_key_mem_340_;
   wire FE_PHN1619_key_mem_355_;
   wire FE_PHN1618_key_mem_365_;
   wire FE_PHN1617_n2133;
   wire FE_PHN1616_key_mem_293_;
   wire FE_PHN1615_key_mem_643_;
   wire FE_PHN1614_key_mem_350_;
   wire FE_PHN1613_key_mem_751_;
   wire FE_PHN1612_n2058;
   wire FE_PHN1611_n1580;
   wire FE_PHN1610_n1908;
   wire FE_PHN1609_key_mem_711_;
   wire FE_PHN1608_n2170;
   wire FE_PHN1607_key_mem_364_;
   wire FE_PHN1606_key_mem_741_;
   wire FE_PHN1605_key_mem_369_;
   wire FE_PHN1604_n1660;
   wire FE_PHN1603_key_mem_330_;
   wire FE_PHN1602_key_mem_765_;
   wire FE_PHN1601_key_mem_294_;
   wire FE_PHN1600_key_mem_303_;
   wire FE_PHN1599_n2171;
   wire FE_PHN1598_key_mem_375_;
   wire FE_PHN1597_n1750;
   wire FE_PHN1596_key_mem_735_;
   wire FE_PHN1595_key_mem_361_;
   wire FE_PHN1594_key_mem_362_;
   wire FE_PHN1593_key_mem_686_;
   wire FE_PHN1592_n1657;
   wire FE_PHN1591_n2064;
   wire FE_PHN1590_key_mem_752_;
   wire FE_PHN1589_key_mem_378_;
   wire FE_PHN1588_key_mem_655_;
   wire FE_PHN1587_key_mem_733_;
   wire FE_PHN1586_key_mem_298_;
   wire FE_PHN1585_n1593;
   wire FE_PHN1584_key_mem_313_;
   wire FE_PHN1583_key_mem_357_;
   wire FE_PHN1582_n1545;
   wire FE_PHN1581_key_mem_672_;
   wire FE_PHN1580_key_mem_372_;
   wire FE_PHN1579_key_mem_678_;
   wire FE_PHN1578_n1418;
   wire FE_PHN1577_key_mem_654_;
   wire FE_PHN1576_n1546;
   wire FE_PHN1575_key_mem_683_;
   wire FE_PHN1574_key_mem_705_;
   wire FE_PHN1573_key_mem_290_;
   wire FE_PHN1572_key_mem_347_;
   wire FE_PHN1571_key_mem_268_;
   wire FE_PHN1570_n1577;
   wire FE_PHN1569_key_mem_670_;
   wire FE_PHN1568_key_mem_720_;
   wire FE_PHN1567_n2057;
   wire FE_PHN1566_n2264;
   wire FE_PHN1565_key_mem_679_;
   wire FE_PHN1564_key_mem_681_;
   wire FE_PHN1563_key_mem_368_;
   wire FE_PHN1562_key_mem_296_;
   wire FE_PHN1561_key_mem_706_;
   wire FE_PHN1560_key_mem_811_;
   wire FE_PHN1559_key_mem_306_;
   wire FE_PHN1558_n2265;
   wire FE_PHN1557_key_mem_305_;
   wire FE_PHN1556_key_mem_725_;
   wire FE_PHN1555_key_mem_320_;
   wire FE_PHN1554_key_mem_282_;
   wire FE_PHN1553_key_mem_257_;
   wire FE_PHN1552_key_mem_763_;
   wire FE_PHN1551_n1739;
   wire FE_PHN1550_key_mem_744_;
   wire FE_PHN1549_key_mem_356_;
   wire FE_PHN1548_n2187;
   wire FE_PHN1547_key_mem_310_;
   wire FE_PHN1546_key_mem_259_;
   wire FE_PHN1545_key_mem_299_;
   wire FE_PHN1544_key_mem_300_;
   wire FE_PHN1543_key_mem_327_;
   wire FE_PHN1542_key_mem_273_;
   wire FE_PHN1541_n1447;
   wire FE_PHN1540_n1419;
   wire FE_PHN1539_n1800;
   wire FE_PHN1538_key_mem_366_;
   wire FE_PHN1537_key_mem_312_;
   wire FE_PHN1536_key_mem_754_;
   wire FE_PHN1535_key_mem_699_;
   wire FE_PHN1534_n1659;
   wire FE_PHN1533_key_mem_337_;
   wire FE_PHN1532_key_mem_806_;
   wire FE_PHN1531_key_mem_762_;
   wire FE_PHN1530_key_mem_719_;
   wire FE_PHN1529_key_mem_314_;
   wire FE_PHN1528_key_mem_729_;
   wire FE_PHN1527_n2183;
   wire FE_PHN1526_n2281;
   wire FE_PHN1525_key_mem_292_;
   wire FE_PHN1524_key_mem_712_;
   wire FE_PHN1523_key_mem_717_;
   wire FE_PHN1522_key_mem_276_;
   wire FE_PHN1521_key_mem_718_;
   wire FE_PHN1520_key_mem_736_;
   wire FE_PHN1519_key_mem_722_;
   wire FE_PHN1518_key_mem_283_;
   wire FE_PHN1517_key_mem_383_;
   wire FE_PHN1516_key_mem_702_;
   wire FE_PHN1515_key_mem_377_;
   wire FE_PHN1514_key_mem_332_;
   wire FE_PHN1513_n2048;
   wire FE_PHN1512_key_mem_664_;
   wire FE_PHN1511_key_mem_295_;
   wire FE_PHN1510_n1738;
   wire FE_PHN1509_n2147;
   wire FE_PHN1508_n1413;
   wire FE_PHN1507_key_mem_304_;
   wire FE_PHN1506_key_mem_690_;
   wire FE_PHN1505_key_mem_658_;
   wire FE_PHN1504_key_mem_271_;
   wire FE_PHN1503_key_mem_382_;
   wire FE_PHN1502_key_mem_642_;
   wire FE_PHN1501_key_mem_381_;
   wire FE_PHN1500_key_mem_749_;
   wire FE_PHN1499_n2107;
   wire FE_PHN1498_key_mem_373_;
   wire FE_PHN1497_n2042;
   wire FE_PHN1496_key_mem_319_;
   wire FE_PHN1495_key_mem_714_;
   wire FE_PHN1494_key_mem_335_;
   wire FE_PHN1493_key_mem_336_;
   wire FE_PHN1492_key_mem_289_;
   wire FE_PHN1491_key_mem_840_;
   wire FE_PHN1490_n2076;
   wire FE_PHN1489_n2263;
   wire FE_PHN1488_n2144;
   wire FE_PHN1487_n1667;
   wire FE_PHN1486_n1752;
   wire FE_PHN1485_n2063;
   wire FE_PHN1484_key_mem_277_;
   wire FE_PHN1483_key_mem_700_;
   wire FE_PHN1482_key_mem_284_;
   wire FE_PHN1481_key_mem_649_;
   wire FE_PHN1480_n1902;
   wire FE_PHN1479_key_mem_326_;
   wire FE_PHN1478_n2106;
   wire FE_PHN1477_key_mem_286_;
   wire FE_PHN1476_key_mem_691_;
   wire FE_PHN1475_key_mem_331_;
   wire FE_PHN1474_n1737;
   wire FE_PHN1473_key_mem_748_;
   wire FE_PHN1472_key_mem_333_;
   wire FE_PHN1471_n2056;
   wire FE_PHN1470_n2050;
   wire FE_PHN1469_key_mem_835_;
   wire FE_PHN1468_n2266;
   wire FE_PHN1467_n1658;
   wire FE_PHN1466_n2124;
   wire FE_PHN1464_key_mem_339_;
   wire FE_PHN1463_n2399;
   wire FE_PHN1446_prev_key1_reg_68_;
   wire FE_PHN1445_prev_key1_reg_69_;
   wire FE_PHN1444_prev_key1_reg_67_;
   wire FE_PHN1442_prev_key1_reg_66_;
   wire FE_PHN1441_prev_key1_reg_64_;
   wire FE_PHN1434_prev_key1_reg_127_;
   wire FE_PHN1429_prev_key1_reg_76_;
   wire FE_PHN1425_prev_key1_reg_81_;
   wire FE_PHN1421_prev_key1_reg_124_;
   wire FE_PHN1416_prev_key1_reg_120_;
   wire FE_PHN1415_prev_key1_reg_75_;
   wire FE_PHN1414_prev_key1_reg_80_;
   wire FE_PHN1413_prev_key1_reg_123_;
   wire FE_PHN1412_prev_key1_reg_85_;
   wire FE_PHN1408_prev_key1_reg_74_;
   wire FE_PHN1406_prev_key1_reg_71_;
   wire FE_PHN1405_prev_key1_reg_82_;
   wire FE_PHN1404_prev_key1_reg_72_;
   wire FE_PHN1402_prev_key1_reg_78_;
   wire FE_PHN1401_prev_key1_reg_73_;
   wire FE_PHN1397_prev_key1_reg_77_;
   wire FE_PHN1395_prev_key1_reg_121_;
   wire FE_PHN1394_prev_key1_reg_65_;
   wire FE_PHN1393_prev_key1_reg_79_;
   wire FE_PHN1392_prev_key1_reg_122_;
   wire FE_PHN1391_prev_key1_reg_125_;
   wire FE_PHN1388_prev_key1_reg_83_;
   wire FE_PHN1375_prev_key1_reg_84_;
   wire FE_PHN1333_n1283;
   wire FE_PHN1326_n1227;
   wire FE_PHN1324_n1029;
   wire FE_PHN1323_n1163;
   wire FE_PHN1322_n1030;
   wire FE_PHN1321_n971;
   wire FE_PHN1318_n972;
   wire FE_PHN1315_n2373;
   wire FE_PHN1314_prev_key1_reg_119_;
   wire FE_PHN1313_prev_key1_reg_118_;
   wire FE_PHN1312_n2381;
   wire FE_PHN1311_n1967;
   wire FE_PHN1263_rcon_reg_1_;
   wire FE_PHN1257_rcon_reg_4_;
   wire FE_PHN1256_prev_key1_reg_112_;
   wire FE_PHN1252_prev_key1_reg_105_;
   wire FE_PHN1251_prev_key1_reg_108_;
   wire FE_PHN1249_prev_key1_reg_116_;
   wire FE_PHN1246_n1736;
   wire FE_PHN1245_prev_key1_reg_99_;
   wire FE_PHN1244_prev_key1_reg_115_;
   wire FE_PHN1241_rcon_reg_5_;
   wire FE_PHN1239_prev_key1_reg_97_;
   wire FE_PHN1238_prev_key1_reg_98_;
   wire FE_PHN1236_prev_key1_reg_113_;
   wire FE_PHN1235_prev_key1_reg_117_;
   wire FE_PHN1234_prev_key1_reg_109_;
   wire FE_PHN1233_prev_key1_reg_106_;
   wire FE_PHN1232_prev_key1_reg_107_;
   wire FE_PHN1231_prev_key1_reg_96_;
   wire FE_PHN1230_prev_key1_reg_53_;
   wire FE_PHN1229_prev_key1_reg_101_;
   wire FE_PHN1227_n2279;
   wire FE_PHN1226_prev_key1_reg_114_;
   wire FE_PHN1225_prev_key1_reg_100_;
   wire FE_PHN1224_prev_key1_reg_103_;
   wire FE_PHN1223_prev_key1_reg_104_;
   wire FE_PHN1221_prev_key1_reg_111_;
   wire FE_PHN1220_prev_key1_reg_102_;
   wire FE_PHN1219_prev_key1_reg_110_;
   wire FE_PHN1211_n2294;
   wire FE_PHN1164_n1282;
   wire FE_PHN1100_n1288;
   wire FE_PHN1098_n1170;
   wire FE_PHN1096_n1022;
   wire FE_PHN1093_n1153;
   wire FE_PHN1092_n1296;
   wire FE_PHN1088_n1295;
   wire FE_PHN1087_prev_key1_reg_44_;
   wire FE_PHN1086_n1166;
   wire FE_PHN1085_n1041;
   wire FE_PHN1084_n1013;
   wire FE_PHN1083_key_mem_1189_;
   wire FE_PHN1081_n1299;
   wire FE_PHN1080_n1280;
   wire FE_PHN1079_prev_key1_reg_32_;
   wire FE_PHN1077_n991;
   wire FE_PHN1076_n1023;
   wire FE_PHN1075_n1290;
   wire FE_PHN1074_prev_key1_reg_50_;
   wire FE_PHN1067_prev_key1_reg_49_;
   wire FE_PHN1066_n908;
   wire FE_PHN1064_prev_key1_reg_45_;
   wire FE_PHN1063_prev_key1_reg_35_;
   wire FE_PHN1062_prev_key1_reg_47_;
   wire FE_PHN1060_prev_key1_reg_33_;
   wire FE_PHN1058_prev_key1_reg_41_;
   wire FE_PHN1057_prev_key1_reg_55_;
   wire FE_PHN1056_prev_key1_reg_37_;
   wire FE_PHN1055_prev_key1_reg_38_;
   wire FE_PHN1054_prev_key1_reg_42_;
   wire FE_PHN1053_prev_key1_reg_36_;
   wire FE_PHN1052_prev_key1_reg_51_;
   wire FE_PHN1051_prev_key1_reg_40_;
   wire FE_PHN1050_prev_key1_reg_54_;
   wire FE_PHN1049_prev_key1_reg_39_;
   wire FE_PHN1048_prev_key1_reg_43_;
   wire FE_PHN1046_n2061;
   wire FE_PHN1045_n1782;
   wire FE_PHN1044_prev_key1_reg_34_;
   wire FE_PHN1043_prev_key1_reg_52_;
   wire FE_PHN1041_n1808;
   wire FE_PHN1040_n1766;
   wire FE_PHN1038_n2418;
   wire FE_PHN1037_n2432;
   wire FE_PHN1036_rcon_reg_3_;
   wire FE_PHN1035_n2350;
   wire FE_PHN1034_rcon_reg_0_;
   wire FE_PHN1033_rcon_reg_2_;
   wire FE_PHN1032_n2868;
   wire FE_PHN1029_key_mem_1193_;
   wire FE_PHN1024_key_mem_1205_;
   wire FE_PHN1023_key_mem_1155_;
   wire FE_PHN1022_n1268;
   wire FE_PHN1021_key_mem_1206_;
   wire FE_PHN1016_n1201;
   wire FE_PHN1015_key_mem_1186_;
   wire FE_PHN1014_key_mem_1253_;
   wire FE_PHN1011_n1076;
   wire FE_PHN1010_key_mem_1222_;
   wire FE_PHN1009_key_mem_1259_;
   wire FE_PHN1008_key_mem_1199_;
   wire FE_PHN1006_key_mem_1219_;
   wire FE_PHN1005_key_mem_1192_;
   wire FE_PHN1000_key_mem_1174_;
   wire FE_PHN999_n1182;
   wire FE_PHN998_n1376;
   wire FE_PHN997_n1386;
   wire FE_PHN996_n1265;
   wire FE_PHN995_n1320;
   wire FE_PHN994_n888;
   wire FE_PHN993_n1379;
   wire FE_PHN992_key_mem_1202_;
   wire FE_PHN991_n1306;
   wire FE_PHN990_key_mem_1270_;
   wire FE_PHN989_key_mem_1157_;
   wire FE_PHN988_n1391;
   wire FE_PHN986_n1121;
   wire FE_PHN984_key_mem_1271_;
   wire FE_PHN983_n1331;
   wire FE_PHN982_n1017;
   wire FE_PHN981_key_mem_1261_;
   wire FE_PHN980_key_mem_1158_;
   wire FE_PHN979_prev_key1_reg_88_;
   wire FE_PHN977_key_mem_1220_;
   wire FE_PHN976_n892;
   wire FE_PHN975_key_mem_1227_;
   wire FE_PHN974_key_mem_1163_;
   wire FE_PHN973_n1196;
   wire FE_PHN972_key_mem_1235_;
   wire FE_PHN971_n1012;
   wire FE_PHN970_n1055;
   wire FE_PHN969_key_mem_1344_;
   wire FE_PHN968_key_mem_1236_;
   wire FE_PHN966_n1385;
   wire FE_PHN965_key_mem_1266_;
   wire FE_PHN964_n1688;
   wire FE_PHN963_n1124;
   wire FE_PHN962_n1184;
   wire FE_PHN961_n1143;
   wire FE_PHN960_key_mem_1228_;
   wire FE_PHN959_n1254;
   wire FE_PHN958_key_mem_1201_;
   wire FE_PHN957_n1396;
   wire FE_PHN956_n1128;
   wire FE_PHN955_key_mem_1198_;
   wire FE_PHN954_key_mem_1063_;
   wire FE_PHN953_key_mem_1200_;
   wire FE_PHN950_n891;
   wire FE_PHN949_key_mem_1231_;
   wire FE_PHN948_n1395;
   wire FE_PHN947_key_mem_1260_;
   wire FE_PHN945_n1185;
   wire FE_PHN944_n1127;
   wire FE_PHN943_key_mem_1195_;
   wire FE_PHN942_key_mem_1203_;
   wire FE_PHN940_prev_key1_reg_95_;
   wire FE_PHN939_key_mem_695_;
   wire FE_PHN938_n944;
   wire FE_PHN937_n990;
   wire FE_PHN936_key_mem_1238_;
   wire FE_PHN935_key_mem_1268_;
   wire FE_PHN934_key_mem_1229_;
   wire FE_PHN933_prev_key1_reg_94_;
   wire FE_PHN932_key_mem_1379_;
   wire FE_PHN930_n946;
   wire FE_PHN929_key_mem_1196_;
   wire FE_PHN928_n994;
   wire FE_PHN924_prev_key1_reg_90_;
   wire FE_PHN923_n1071;
   wire FE_PHN922_prev_key1_reg_89_;
   wire FE_PHN921_prev_key1_reg_91_;
   wire FE_PHN919_prev_key1_reg_92_;
   wire FE_PHN917_key_mem_676_;
   wire FE_PHN916_n1600;
   wire FE_PHN915_key_mem_371_;
   wire FE_PHN914_key_mem_652_;
   wire FE_PHN913_n2157;
   wire FE_PHN912_rcon_reg_7_;
   wire FE_PHN896_prev_key1_reg_61_;
   wire FE_PHN827_n2122;
   wire FE_PHN819_key_mem_1176_;
   wire FE_PHN817_key_mem_1240_;
   wire FE_PHN812_n1206;
   wire FE_PHN811_key_mem_1247_;
   wire FE_PHN810_n1059;
   wire FE_PHN808_key_mem_1182_;
   wire FE_PHN807_n1146;
   wire FE_PHN806_n1317;
   wire FE_PHN803_n1190;
   wire FE_PHN802_key_mem_1273_;
   wire FE_PHN800_key_mem_1214_;
   wire FE_PHN798_key_mem_1166_;
   wire FE_PHN797_key_mem_1212_;
   wire FE_PHN796_n1342;
   wire FE_PHN794_key_mem_1246_;
   wire FE_PHN792_key_mem_1277_;
   wire FE_PHN791_key_mem_1177_;
   wire FE_PHN789_n1205;
   wire FE_PHN788_key_mem_1372_;
   wire FE_PHN786_key_mem_1208_;
   wire FE_PHN785_key_mem_1218_;
   wire FE_PHN783_key_mem_1209_;
   wire FE_PHN782_key_mem_1213_;
   wire FE_PHN780_key_mem_1276_;
   wire FE_PHN779_key_mem_1249_;
   wire FE_PHN777_key_mem_1234_;
   wire FE_PHN776_key_mem_1239_;
   wire FE_PHN775_key_mem_1156_;
   wire FE_PHN774_key_mem_1345_;
   wire FE_PHN773_key_mem_1245_;
   wire FE_PHN772_key_mem_760_;
   wire FE_PHN771_key_mem_1243_;
   wire FE_PHN770_key_mem_1241_;
   wire FE_PHN769_n1323;
   wire FE_PHN768_key_mem_1173_;
   wire FE_PHN767_key_mem_1242_;
   wire FE_PHN766_key_mem_1274_;
   wire FE_PHN765_key_mem_1211_;
   wire FE_PHN764_key_mem_287_;
   wire FE_PHN763_key_mem_275_;
   wire FE_PHN762_key_mem_767_;
   wire FE_PHN760_key_mem_1179_;
   wire FE_PHN758_key_mem_703_;
   wire FE_PHN757_prev_key1_reg_93_;
   wire FE_PHN756_key_mem_766_;
   wire FE_PHN755_key_mem_379_;
   wire FE_PHN754_key_mem_657_;
   wire FE_PHN748_keymem_sboxw_6_;
   wire FE_PHN747_n2364;
   wire FE_PHN746_prev_key1_reg_58_;
   wire FE_PHN745_prev_key1_reg_59_;
   wire FE_PHN744_prev_key1_reg_57_;
   wire FE_PHN743_prev_key1_reg_63_;
   wire FE_PHN741_prev_key1_reg_60_;
   wire FE_PHN740_prev_key1_reg_62_;
   wire FE_PHN739_n1244;
   wire FE_PHN738_n1365;
   wire FE_PHN737_n1354;
   wire FE_PHN736_n1219;
   wire FE_PHN735_n1225;
   wire FE_PHN734_n1345;
   wire FE_PHN733_n1360;
   wire FE_PHN732_n1343;
   wire FE_PHN731_n953;
   wire FE_PHN730_n1112;
   wire FE_PHN728_n1236;
   wire FE_PHN727_n968;
   wire FE_PHN726_n1095;
   wire FE_PHN724_n1107;
   wire FE_PHN723_n1366;
   wire FE_PHN722_n1335;
   wire FE_PHN721_n1111;
   wire FE_PHN720_n1088;
   wire FE_PHN719_n978;
   wire FE_PHN718_n962;
   wire FE_PHN717_n987;
   wire FE_PHN716_n1105;
   wire FE_PHN715_n2372;
   wire FE_PHN714_n2374;
   wire FE_PHN713_n1114;
   wire FE_PHN712_n955;
   wire FE_PHN710_n1364;
   wire FE_PHN709_n985;
   wire FE_PHN708_n975;
   wire FE_PHN707_n1336;
   wire FE_PHN706_n1102;
   wire FE_PHN705_n629;
   wire FE_PHN700_key_mem_1265_;
   wire FE_PHN699_key_mem_1254_;
   wire FE_PHN698_key_mem_1172_;
   wire FE_PHN696_key_mem_1194_;
   wire FE_PHN694_key_mem_1232_;
   wire FE_PHN692_key_mem_1226_;
   wire FE_PHN691_key_mem_1248_;
   wire FE_PHN689_key_mem_1223_;
   wire FE_PHN688_key_mem_1252_;
   wire FE_PHN686_key_mem_1250_;
   wire FE_PHN684_key_mem_640_;
   wire FE_PHN683_key_mem_641_;
   wire FE_PHN646_n1308;
   wire FE_PHN638_n1048;
   wire FE_PHN635_n1373;
   wire FE_PHN633_n1305;
   wire FE_PHN632_n1175;
   wire FE_PHN631_n917;
   wire FE_PHN628_n923;
   wire FE_PHN627_n1768;
   wire FE_PHN626_n1439;
   wire FE_PHN625_n649;
   wire FE_PHN624_n551;
   wire FE_PHN623_n544;
   wire FE_PHN622_n543;
   wire FE_PHN621_n561;
   wire FE_PHN620_n554;
   wire FE_PHN619_n555;
   wire FE_PHN618_n562;
   wire FE_PHN617_n570;
   wire FE_PHN616_n553;
   wire FE_PHN615_n563;
   wire FE_PHN614_n556;
   wire FE_PHN613_n569;
   wire FE_PHN612_n572;
   wire FE_PHN611_n567;
   wire FE_PHN610_n573;
   wire FE_PHN609_n574;
   wire FE_PHN608_n564;
   wire FE_PHN607_n566;
   wire FE_PHN606_n571;
   wire FE_PHN605_n568;
   wire FE_PHN594_key_mem_1225_;
   wire FE_PHN593_n1381;
   wire FE_PHN592_key_mem_1390_;
   wire FE_PHN591_key_mem_1230_;
   wire FE_PHN590_n1389;
   wire FE_PHN589_n1082;
   wire FE_PHN588_n1259;
   wire FE_PHN587_key_mem_1161_;
   wire FE_PHN586_n1132;
   wire FE_PHN585_key_mem_1175_;
   wire FE_PHN584_key_mem_1159_;
   wire FE_PHN583_key_mem_1257_;
   wire FE_PHN582_key_mem_1170_;
   wire FE_PHN581_n1004;
   wire FE_PHN580_key_mem_743_;
   wire FE_PHN579_n650;
   wire FE_PHN578_n600;
   wire FE_PHN577_n593;
   wire FE_PHN576_n584;
   wire FE_PHN575_n594;
   wire FE_PHN574_n583;
   wire FE_PHN573_n654;
   wire FE_PHN572_n664;
   wire FE_PHN571_n656;
   wire FE_PHN570_n653;
   wire FE_PHN569_n651;
   wire FE_PHN568_n550;
   wire FE_PHN567_n549;
   wire FE_PHN566_n665;
   wire FE_PHN565_n596;
   wire FE_PHN564_n648;
   wire FE_PHN563_n667;
   wire FE_PHN562_n666;
   wire FE_PHN561_n601;
   wire FE_PHN560_n658;
   wire FE_PHN559_n598;
   wire FE_PHN558_n652;
   wire FE_PHN557_n602;
   wire FE_PHN556_n595;
   wire FE_PHN555_n605;
   wire FE_PHN554_n659;
   wire FE_PHN553_n670;
   wire FE_PHN552_n657;
   wire FE_PHN551_n545;
   wire FE_PHN550_n668;
   wire FE_PHN549_n587;
   wire FE_PHN548_n546;
   wire FE_PHN547_n580;
   wire FE_PHN546_n603;
   wire FE_PHN545_n599;
   wire FE_PHN544_n547;
   wire FE_PHN543_n588;
   wire FE_PHN542_n586;
   wire FE_PHN541_n660;
   wire FE_PHN540_n606;
   wire FE_PHN539_n585;
   wire FE_PHN538_n604;
   wire FE_PHN537_n669;
   wire FE_PHN432_key_mem_1256_;
   wire FE_PHN431_key_mem_1224_;
   wire FE_PHN430_key_mem_1167_;
   wire FE_PHN429_key_mem_1162_;
   wire FE_PHN428_n1161;
   wire FE_PHN427_key_mem_1258_;
   wire FE_PHN426_key_mem_1184_;
   wire FE_PHN425_key_mem_1264_;
   wire FE_PHN424_key_mem_367_;
   wire FE_PHN423_n607;
   wire FE_PHN422_n608;
   wire FE_PHN421_n590;
   wire FE_PHN420_n592;
   wire FE_PHN419_n589;
   wire FE_PHN418_n548;
   wire FE_PHN417_n591;
   wire FE_PHN416_n597;
   wire FE_PHN411_n6;
   wire FE_PHN409_n624;
   wire FE_PHN408_n640;
   wire FE_PHN407_n645;
   wire FE_PHN406_n646;
   wire FE_PHN405_n613;
   wire FE_PHN404_n614;
   wire FE_PHN403_n622;
   wire FE_PHN402_n621;
   wire FE_PHN401_n639;
   wire FE_PHN400_n641;
   wire FE_PHN399_n643;
   wire FE_PHN398_n627;
   wire FE_PHN397_n642;
   wire FE_PHN396_n632;
   wire FE_PHN395_n644;
   wire FE_PHN394_n634;
   wire FE_PHN393_n609;
   wire FE_PHN392_n610;
   wire FE_PHN391_n633;
   wire FE_PHN390_n628;
   wire FE_PHN389_n618;
   wire FE_PHN388_n626;
   wire FE_PHN387_n625;
   wire FE_PHN386_n611;
   wire FE_PHN385_n617;
   wire FE_PHN384_n620;
   wire FE_PHN383_n638;
   wire FE_PHN382_n619;
   wire FE_PHN381_n636;
   wire FE_PHN380_n637;
   wire FE_PHN379_n635;
   wire FE_PHN360_prev_key1_reg_86_;
   wire FE_PHN359_prev_key1_reg_87_;
   wire FE_PHN357_key_mem_1154_;
   wire FE_PHN349_n581;
   wire FE_PHN348_n647;
   wire FE_PHN347_n582;
   wire FE_PHN346_n579;
   wire FE_PHN345_n578;
   wire FE_PHN344_n576;
   wire FE_PHN343_n577;
   wire FE_PHN342_n575;
   wire FE_PHN327_n655;
   wire FE_PHN326_n612;
   wire FE_PHN325_n662;
   wire FE_PHN324_n663;
   wire FE_PHN323_n661;
   wire FE_PHN290_key_mem_ctrl_reg_0_;
   wire FE_PHN283_n2433;
   wire FE_PHN265_keymem_sboxw_7_;
   wire FE_PHN254_n689;
   wire FE_PHN198_round_ctr_reg_0_;
   wire FE_PHN178_round_ctr_reg_2_;
   wire FE_PHN155_n3;
   wire FE_PHN120_key_mem_ctrl_reg_1_;
   wire FE_PHN116_round_ctr_reg_3_;
   wire FE_PHN112_round_ctr_reg_1_;
   wire FE_OFN109_n23;
   wire FE_OFN108_n21;
   wire FE_OFN107_n21;
   wire FE_OFN106_n22;
   wire FE_OFN105_n2763;
   wire FE_OFN104_n27;
   wire FE_OFN103_n27;
   wire FE_OFN102_n31;
   wire FE_OFN101_n30;
   wire FE_OFN100_n2800;
   wire FE_OFN99_n2811;
   wire FE_OFN96_n674;
   wire FE_OFN95_n674;
   wire FE_OFN94_n674;
   wire FE_OFN93_n674;
   wire FE_OFN92_n674;
   wire FE_OFN91_n690;
   wire FE_OFN90_n690;
   wire FE_OFN89_n1;
   wire FE_OFN88_n1;
   wire FE_OFN87_n1;
   wire FE_OFN86_n1;
   wire FE_OFN85_n1;
   wire FE_OFN84_n1;
   wire FE_OFN83_n672;
   wire FE_OFN82_n672;
   wire FE_OFN81_n672;
   wire FE_OFN80_n672;
   wire FE_OFN79_n672;
   wire FE_OFN78_n676;
   wire FE_OFN77_n676;
   wire FE_OFN76_n676;
   wire FE_OFN57_reset_n;
   wire FE_OFN41_reset_n;
   wire FE_OFN36_reset_n;
   wire FE_OFN33_n683;
   wire FE_OFN32_n683;
   wire FE_OFN31_n683;
   wire FE_OFN30_n687;
   wire FE_OFN29_n687;
   wire FE_OFN28_n687;
   wire FE_OFN27_n685;
   wire FE_OFN26_n685;
   wire FE_OFN25_n685;
   wire FE_OFN24_n685;
   wire FE_OFN23_n681;
   wire FE_OFN22_n681;
   wire FE_OFN21_n681;
   wire FE_OFN20_n681;
   wire FE_OFN19_n681;
   wire FE_OFN18_n678;
   wire FE_OFN17_n678;
   wire FE_OFN16_n678;
   wire FE_OFN15_n678;
   wire FE_OFN14_n688;
   wire FE_OFN13_n688;
   wire FE_OFN12_n688;
   wire FE_OFN11_n688;
   wire FE_OFN10_n688;
   wire FE_OFN9_n684;
   wire FE_OFN8_n684;
   wire FE_OFN7_n684;
   wire FE_OFN6_n684;
   wire FE_OFN5_n682;
   wire FE_OFN4_n682;
   wire FE_OFN3_n682;
   wire FE_OFN2_n682;
   wire FE_OFN1_n682;
   wire n6;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n27;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire n478;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire n556;
   wire n557;
   wire n558;
   wire n559;
   wire n560;
   wire n561;
   wire n562;
   wire n563;
   wire n564;
   wire n565;
   wire n566;
   wire n567;
   wire n568;
   wire n569;
   wire n570;
   wire n571;
   wire n572;
   wire n573;
   wire n574;
   wire n575;
   wire n576;
   wire n577;
   wire n578;
   wire n579;
   wire n580;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire n593;
   wire n594;
   wire n595;
   wire n596;
   wire n597;
   wire n598;
   wire n599;
   wire n600;
   wire n601;
   wire n602;
   wire n603;
   wire n604;
   wire n605;
   wire n606;
   wire n607;
   wire n608;
   wire n609;
   wire n610;
   wire n611;
   wire n612;
   wire n613;
   wire n614;
   wire n615;
   wire n616;
   wire n617;
   wire n618;
   wire n619;
   wire n620;
   wire n621;
   wire n622;
   wire n623;
   wire n624;
   wire n625;
   wire n626;
   wire n627;
   wire n628;
   wire n629;
   wire n630;
   wire n631;
   wire n632;
   wire n633;
   wire n634;
   wire n635;
   wire n636;
   wire n637;
   wire n638;
   wire n639;
   wire n640;
   wire n641;
   wire n642;
   wire n643;
   wire n644;
   wire n645;
   wire n646;
   wire n647;
   wire n648;
   wire n649;
   wire n650;
   wire n651;
   wire n652;
   wire n653;
   wire n654;
   wire n655;
   wire n656;
   wire n657;
   wire n658;
   wire n659;
   wire n660;
   wire n661;
   wire n662;
   wire n663;
   wire n664;
   wire n665;
   wire n666;
   wire n667;
   wire n668;
   wire n669;
   wire n670;
   wire n672;
   wire n673;
   wire n674;
   wire n675;
   wire n676;
   wire n677;
   wire n678;
   wire n679;
   wire n680;
   wire n681;
   wire n682;
   wire n683;
   wire n684;
   wire n685;
   wire n686;
   wire n687;
   wire n688;
   wire n689;
   wire n690;
   wire n691;
   wire n692;
   wire n693;
   wire n694;
   wire n695;
   wire n696;
   wire n697;
   wire n698;
   wire n699;
   wire n700;
   wire n701;
   wire n702;
   wire n703;
   wire n704;
   wire n705;
   wire n706;
   wire n707;
   wire n708;
   wire n709;
   wire n710;
   wire n711;
   wire n712;
   wire n713;
   wire n714;
   wire n715;
   wire n716;
   wire n717;
   wire n718;
   wire n719;
   wire n720;
   wire n721;
   wire n722;
   wire n723;
   wire n724;
   wire n725;
   wire n726;
   wire n727;
   wire n728;
   wire n729;
   wire n730;
   wire n731;
   wire n732;
   wire n733;
   wire n734;
   wire n735;
   wire n736;
   wire n737;
   wire n738;
   wire n739;
   wire n740;
   wire n741;
   wire n742;
   wire n743;
   wire n744;
   wire n745;
   wire n746;
   wire n747;
   wire n748;
   wire n749;
   wire n750;
   wire n751;
   wire n752;
   wire n753;
   wire n754;
   wire n755;
   wire n756;
   wire n757;
   wire n758;
   wire n759;
   wire n760;
   wire n761;
   wire n762;
   wire n763;
   wire n764;
   wire n765;
   wire n766;
   wire n767;
   wire n768;
   wire n769;
   wire n770;
   wire n771;
   wire n772;
   wire n773;
   wire n774;
   wire n775;
   wire n776;
   wire n777;
   wire n778;
   wire n779;
   wire n780;
   wire n781;
   wire n782;
   wire n783;
   wire n784;
   wire n785;
   wire n786;
   wire n787;
   wire n788;
   wire n789;
   wire n790;
   wire n791;
   wire n792;
   wire n793;
   wire n794;
   wire n795;
   wire n796;
   wire n797;
   wire n798;
   wire n799;
   wire n800;
   wire n801;
   wire n802;
   wire n803;
   wire n804;
   wire n805;
   wire n806;
   wire n807;
   wire n808;
   wire n809;
   wire n810;
   wire n811;
   wire n812;
   wire n813;
   wire n814;
   wire n815;
   wire n816;
   wire n817;
   wire n818;
   wire n819;
   wire n820;
   wire n821;
   wire n822;
   wire n823;
   wire n824;
   wire n825;
   wire n826;
   wire n827;
   wire n828;
   wire n829;
   wire n830;
   wire n831;
   wire n832;
   wire n833;
   wire n834;
   wire n835;
   wire n836;
   wire n837;
   wire n838;
   wire n839;
   wire n840;
   wire n841;
   wire n842;
   wire n843;
   wire n844;
   wire n845;
   wire n846;
   wire n847;
   wire n848;
   wire n849;
   wire n850;
   wire n851;
   wire n852;
   wire n853;
   wire n854;
   wire n855;
   wire n856;
   wire n857;
   wire n858;
   wire n859;
   wire n860;
   wire n861;
   wire n862;
   wire n863;
   wire n864;
   wire n865;
   wire n866;
   wire n867;
   wire n868;
   wire n869;
   wire n870;
   wire n871;
   wire n872;
   wire n873;
   wire n874;
   wire n875;
   wire n876;
   wire n877;
   wire n878;
   wire n879;
   wire n880;
   wire n881;
   wire n882;
   wire n883;
   wire n884;
   wire n885;
   wire n886;
   wire n887;
   wire n888;
   wire n889;
   wire n890;
   wire n891;
   wire n892;
   wire n893;
   wire n894;
   wire n895;
   wire n896;
   wire n897;
   wire n898;
   wire n899;
   wire n900;
   wire n901;
   wire n902;
   wire n903;
   wire n904;
   wire n905;
   wire n906;
   wire n907;
   wire n908;
   wire n909;
   wire n910;
   wire n911;
   wire n912;
   wire n913;
   wire n914;
   wire n915;
   wire n916;
   wire n917;
   wire n918;
   wire n919;
   wire n920;
   wire n921;
   wire n922;
   wire n923;
   wire n924;
   wire n925;
   wire n926;
   wire n927;
   wire n928;
   wire n929;
   wire n930;
   wire n931;
   wire n932;
   wire n933;
   wire n934;
   wire n935;
   wire n936;
   wire n937;
   wire n938;
   wire n939;
   wire n940;
   wire n941;
   wire n942;
   wire n943;
   wire n944;
   wire n945;
   wire n946;
   wire n947;
   wire n948;
   wire n949;
   wire n950;
   wire n951;
   wire n952;
   wire n953;
   wire n954;
   wire n955;
   wire n956;
   wire n957;
   wire n958;
   wire n959;
   wire n960;
   wire n961;
   wire n962;
   wire n963;
   wire n964;
   wire n965;
   wire n966;
   wire n967;
   wire n968;
   wire n969;
   wire n970;
   wire n971;
   wire n972;
   wire n973;
   wire n974;
   wire n975;
   wire n976;
   wire n977;
   wire n978;
   wire n979;
   wire n980;
   wire n981;
   wire n982;
   wire n983;
   wire n984;
   wire n985;
   wire n986;
   wire n987;
   wire n988;
   wire n989;
   wire n990;
   wire n991;
   wire n992;
   wire n993;
   wire n994;
   wire n995;
   wire n996;
   wire n997;
   wire n998;
   wire n999;
   wire n1000;
   wire n1001;
   wire n1002;
   wire n1003;
   wire n1004;
   wire n1005;
   wire n1006;
   wire n1007;
   wire n1008;
   wire n1009;
   wire n1010;
   wire n1011;
   wire n1012;
   wire n1013;
   wire n1014;
   wire n1015;
   wire n1016;
   wire n1017;
   wire n1018;
   wire n1019;
   wire n1020;
   wire n1021;
   wire n1022;
   wire n1023;
   wire n1024;
   wire n1025;
   wire n1026;
   wire n1027;
   wire n1028;
   wire n1029;
   wire n1030;
   wire n1031;
   wire n1032;
   wire n1033;
   wire n1034;
   wire n1035;
   wire n1036;
   wire n1037;
   wire n1038;
   wire n1039;
   wire n1040;
   wire n1041;
   wire n1042;
   wire n1043;
   wire n1044;
   wire n1045;
   wire n1046;
   wire n1047;
   wire n1048;
   wire n1049;
   wire n1050;
   wire n1051;
   wire n1052;
   wire n1053;
   wire n1054;
   wire n1055;
   wire n1056;
   wire n1057;
   wire n1058;
   wire n1059;
   wire n1060;
   wire n1061;
   wire n1062;
   wire n1063;
   wire n1064;
   wire n1065;
   wire n1066;
   wire n1067;
   wire n1068;
   wire n1069;
   wire n1070;
   wire n1071;
   wire n1072;
   wire n1073;
   wire n1074;
   wire n1075;
   wire n1076;
   wire n1077;
   wire n1078;
   wire n1079;
   wire n1080;
   wire n1081;
   wire n1082;
   wire n1083;
   wire n1084;
   wire n1085;
   wire n1086;
   wire n1087;
   wire n1088;
   wire n1089;
   wire n1090;
   wire n1091;
   wire n1092;
   wire n1093;
   wire n1094;
   wire n1095;
   wire n1096;
   wire n1097;
   wire n1098;
   wire n1099;
   wire n1100;
   wire n1101;
   wire n1102;
   wire n1103;
   wire n1104;
   wire n1105;
   wire n1106;
   wire n1107;
   wire n1108;
   wire n1109;
   wire n1110;
   wire n1111;
   wire n1112;
   wire n1113;
   wire n1114;
   wire n1115;
   wire n1116;
   wire n1117;
   wire n1118;
   wire n1119;
   wire n1120;
   wire n1121;
   wire n1122;
   wire n1123;
   wire n1124;
   wire n1125;
   wire n1126;
   wire n1127;
   wire n1128;
   wire n1129;
   wire n1130;
   wire n1131;
   wire n1132;
   wire n1133;
   wire n1134;
   wire n1135;
   wire n1136;
   wire n1137;
   wire n1138;
   wire n1139;
   wire n1140;
   wire n1141;
   wire n1142;
   wire n1143;
   wire n1144;
   wire n1145;
   wire n1146;
   wire n1147;
   wire n1148;
   wire n1149;
   wire n1150;
   wire n1151;
   wire n1152;
   wire n1153;
   wire n1154;
   wire n1155;
   wire n1156;
   wire n1157;
   wire n1158;
   wire n1159;
   wire n1160;
   wire n1161;
   wire n1162;
   wire n1163;
   wire n1164;
   wire n1165;
   wire n1166;
   wire n1167;
   wire n1168;
   wire n1169;
   wire n1170;
   wire n1171;
   wire n1172;
   wire n1173;
   wire n1174;
   wire n1175;
   wire n1176;
   wire n1177;
   wire n1178;
   wire n1179;
   wire n1180;
   wire n1181;
   wire n1182;
   wire n1183;
   wire n1184;
   wire n1185;
   wire n1186;
   wire n1187;
   wire n1188;
   wire n1189;
   wire n1190;
   wire n1191;
   wire n1192;
   wire n1193;
   wire n1194;
   wire n1195;
   wire n1196;
   wire n1197;
   wire n1198;
   wire n1199;
   wire n1200;
   wire n1201;
   wire n1202;
   wire n1203;
   wire n1204;
   wire n1205;
   wire n1206;
   wire n1207;
   wire n1208;
   wire n1209;
   wire n1210;
   wire n1211;
   wire n1212;
   wire n1213;
   wire n1214;
   wire n1215;
   wire n1216;
   wire n1217;
   wire n1218;
   wire n1219;
   wire n1220;
   wire n1221;
   wire n1222;
   wire n1223;
   wire n1224;
   wire n1225;
   wire n1226;
   wire n1227;
   wire n1228;
   wire n1229;
   wire n1230;
   wire n1231;
   wire n1232;
   wire n1233;
   wire n1234;
   wire n1235;
   wire n1236;
   wire n1237;
   wire n1238;
   wire n1239;
   wire n1240;
   wire n1241;
   wire n1242;
   wire n1243;
   wire n1244;
   wire n1245;
   wire n1246;
   wire n1247;
   wire n1248;
   wire n1249;
   wire n1250;
   wire n1251;
   wire n1252;
   wire n1253;
   wire n1254;
   wire n1255;
   wire n1256;
   wire n1257;
   wire n1258;
   wire n1259;
   wire n1260;
   wire n1261;
   wire n1262;
   wire n1263;
   wire n1264;
   wire n1265;
   wire n1266;
   wire n1267;
   wire n1268;
   wire n1269;
   wire n1270;
   wire n1271;
   wire n1272;
   wire n1273;
   wire n1274;
   wire n1275;
   wire n1276;
   wire n1277;
   wire n1278;
   wire n1279;
   wire n1280;
   wire n1281;
   wire n1282;
   wire n1283;
   wire n1284;
   wire n1285;
   wire n1286;
   wire n1287;
   wire n1288;
   wire n1289;
   wire n1290;
   wire n1291;
   wire n1292;
   wire n1293;
   wire n1294;
   wire n1295;
   wire n1296;
   wire n1297;
   wire n1298;
   wire n1299;
   wire n1300;
   wire n1301;
   wire n1302;
   wire n1303;
   wire n1304;
   wire n1305;
   wire n1306;
   wire n1307;
   wire n1308;
   wire n1309;
   wire n1310;
   wire n1311;
   wire n1312;
   wire n1313;
   wire n1314;
   wire n1315;
   wire n1316;
   wire n1317;
   wire n1318;
   wire n1319;
   wire n1320;
   wire n1321;
   wire n1322;
   wire n1323;
   wire n1324;
   wire n1325;
   wire n1326;
   wire n1327;
   wire n1328;
   wire n1329;
   wire n1330;
   wire n1331;
   wire n1332;
   wire n1333;
   wire n1334;
   wire n1335;
   wire n1336;
   wire n1337;
   wire n1338;
   wire n1339;
   wire n1340;
   wire n1341;
   wire n1342;
   wire n1343;
   wire n1344;
   wire n1345;
   wire n1346;
   wire n1347;
   wire n1348;
   wire n1349;
   wire n1350;
   wire n1351;
   wire n1352;
   wire n1353;
   wire n1354;
   wire n1355;
   wire n1356;
   wire n1357;
   wire n1358;
   wire n1359;
   wire n1360;
   wire n1361;
   wire n1362;
   wire n1363;
   wire n1364;
   wire n1365;
   wire n1366;
   wire n1367;
   wire n1368;
   wire n1369;
   wire n1370;
   wire n1371;
   wire n1372;
   wire n1373;
   wire n1374;
   wire n1375;
   wire n1376;
   wire n1377;
   wire n1378;
   wire n1379;
   wire n1380;
   wire n1381;
   wire n1382;
   wire n1383;
   wire n1384;
   wire n1385;
   wire n1386;
   wire n1387;
   wire n1388;
   wire n1389;
   wire n1390;
   wire n1391;
   wire n1392;
   wire n1393;
   wire n1394;
   wire n1395;
   wire n1396;
   wire n1397;
   wire n1398;
   wire n1399;
   wire n1400;
   wire n1401;
   wire n1402;
   wire n1403;
   wire n1404;
   wire n1405;
   wire n1406;
   wire n1407;
   wire n1408;
   wire n1409;
   wire n1410;
   wire n1411;
   wire n1412;
   wire n1413;
   wire n1414;
   wire n1415;
   wire n1416;
   wire n1417;
   wire n1418;
   wire n1419;
   wire n1420;
   wire n1421;
   wire n1422;
   wire n1423;
   wire n1424;
   wire n1425;
   wire n1426;
   wire n1427;
   wire n1428;
   wire n1429;
   wire n1430;
   wire n1431;
   wire n1432;
   wire n1433;
   wire n1434;
   wire n1435;
   wire n1436;
   wire n1437;
   wire n1438;
   wire n1439;
   wire n1440;
   wire n1441;
   wire n1442;
   wire n1443;
   wire n1444;
   wire n1445;
   wire n1446;
   wire n1447;
   wire n1448;
   wire n1449;
   wire n1450;
   wire n1451;
   wire n1452;
   wire n1453;
   wire n1454;
   wire n1455;
   wire n1456;
   wire n1457;
   wire n1458;
   wire n1459;
   wire n1460;
   wire n1461;
   wire n1462;
   wire n1463;
   wire n1464;
   wire n1465;
   wire n1466;
   wire n1467;
   wire n1468;
   wire n1469;
   wire n1470;
   wire n1471;
   wire n1472;
   wire n1473;
   wire n1474;
   wire n1475;
   wire n1476;
   wire n1477;
   wire n1478;
   wire n1479;
   wire n1480;
   wire n1481;
   wire n1482;
   wire n1483;
   wire n1484;
   wire n1485;
   wire n1486;
   wire n1487;
   wire n1488;
   wire n1489;
   wire n1490;
   wire n1491;
   wire n1492;
   wire n1493;
   wire n1494;
   wire n1495;
   wire n1496;
   wire n1497;
   wire n1498;
   wire n1499;
   wire n1500;
   wire n1501;
   wire n1502;
   wire n1503;
   wire n1504;
   wire n1505;
   wire n1506;
   wire n1507;
   wire n1508;
   wire n1509;
   wire n1510;
   wire n1511;
   wire n1512;
   wire n1513;
   wire n1514;
   wire n1515;
   wire n1516;
   wire n1517;
   wire n1518;
   wire n1519;
   wire n1520;
   wire n1521;
   wire n1522;
   wire n1523;
   wire n1524;
   wire n1525;
   wire n1526;
   wire n1527;
   wire n1528;
   wire n1529;
   wire n1530;
   wire n1531;
   wire n1532;
   wire n1533;
   wire n1534;
   wire n1535;
   wire n1536;
   wire n1537;
   wire n1538;
   wire n1539;
   wire n1540;
   wire n1541;
   wire n1542;
   wire n1543;
   wire n1544;
   wire n1545;
   wire n1546;
   wire n1547;
   wire n1548;
   wire n1549;
   wire n1550;
   wire n1551;
   wire n1552;
   wire n1553;
   wire n1554;
   wire n1555;
   wire n1556;
   wire n1557;
   wire n1558;
   wire n1559;
   wire n1560;
   wire n1561;
   wire n1562;
   wire n1563;
   wire n1564;
   wire n1565;
   wire n1566;
   wire n1567;
   wire n1568;
   wire n1569;
   wire n1570;
   wire n1571;
   wire n1572;
   wire n1573;
   wire n1574;
   wire n1575;
   wire n1576;
   wire n1577;
   wire n1578;
   wire n1579;
   wire n1580;
   wire n1581;
   wire n1582;
   wire n1583;
   wire n1584;
   wire n1585;
   wire n1586;
   wire n1587;
   wire n1588;
   wire n1589;
   wire n1590;
   wire n1591;
   wire n1592;
   wire n1593;
   wire n1594;
   wire n1595;
   wire n1596;
   wire n1597;
   wire n1598;
   wire n1599;
   wire n1600;
   wire n1601;
   wire n1602;
   wire n1603;
   wire n1604;
   wire n1605;
   wire n1606;
   wire n1607;
   wire n1608;
   wire n1609;
   wire n1610;
   wire n1611;
   wire n1612;
   wire n1613;
   wire n1614;
   wire n1615;
   wire n1616;
   wire n1617;
   wire n1618;
   wire n1619;
   wire n1620;
   wire n1621;
   wire n1622;
   wire n1623;
   wire n1624;
   wire n1625;
   wire n1626;
   wire n1627;
   wire n1628;
   wire n1629;
   wire n1630;
   wire n1631;
   wire n1632;
   wire n1633;
   wire n1634;
   wire n1635;
   wire n1636;
   wire n1637;
   wire n1638;
   wire n1639;
   wire n1640;
   wire n1641;
   wire n1642;
   wire n1643;
   wire n1644;
   wire n1645;
   wire n1646;
   wire n1647;
   wire n1648;
   wire n1649;
   wire n1650;
   wire n1651;
   wire n1652;
   wire n1653;
   wire n1654;
   wire n1655;
   wire n1656;
   wire n1657;
   wire n1658;
   wire n1659;
   wire n1660;
   wire n1661;
   wire n1662;
   wire n1663;
   wire n1664;
   wire n1665;
   wire n1666;
   wire n1667;
   wire n1668;
   wire n1669;
   wire n1670;
   wire n1671;
   wire n1672;
   wire n1673;
   wire n1674;
   wire n1675;
   wire n1676;
   wire n1677;
   wire n1678;
   wire n1679;
   wire n1680;
   wire n1681;
   wire n1682;
   wire n1683;
   wire n1684;
   wire n1685;
   wire n1686;
   wire n1687;
   wire n1688;
   wire n1689;
   wire n1690;
   wire n1691;
   wire n1692;
   wire n1693;
   wire n1694;
   wire n1695;
   wire n1696;
   wire n1697;
   wire n1698;
   wire n1699;
   wire n1700;
   wire n1701;
   wire n1702;
   wire n1703;
   wire n1704;
   wire n1705;
   wire n1706;
   wire n1707;
   wire n1708;
   wire n1709;
   wire n1710;
   wire n1711;
   wire n1712;
   wire n1713;
   wire n1714;
   wire n1715;
   wire n1716;
   wire n1717;
   wire n1718;
   wire n1719;
   wire n1720;
   wire n1721;
   wire n1722;
   wire n1723;
   wire n1724;
   wire n1725;
   wire n1726;
   wire n1727;
   wire n1728;
   wire n1729;
   wire n1730;
   wire n1731;
   wire n1732;
   wire n1733;
   wire n1734;
   wire n1735;
   wire n1736;
   wire n1737;
   wire n1738;
   wire n1739;
   wire n1740;
   wire n1741;
   wire n1742;
   wire n1743;
   wire n1744;
   wire n1745;
   wire n1746;
   wire n1747;
   wire n1748;
   wire n1749;
   wire n1750;
   wire n1751;
   wire n1752;
   wire n1753;
   wire n1754;
   wire n1755;
   wire n1756;
   wire n1757;
   wire n1758;
   wire n1759;
   wire n1760;
   wire n1761;
   wire n1762;
   wire n1763;
   wire n1764;
   wire n1765;
   wire n1766;
   wire n1767;
   wire n1768;
   wire n1769;
   wire n1770;
   wire n1771;
   wire n1772;
   wire n1773;
   wire n1774;
   wire n1775;
   wire n1776;
   wire n1777;
   wire n1778;
   wire n1779;
   wire n1780;
   wire n1781;
   wire n1782;
   wire n1783;
   wire n1784;
   wire n1785;
   wire n1786;
   wire n1787;
   wire n1788;
   wire n1789;
   wire n1790;
   wire n1791;
   wire n1792;
   wire n1793;
   wire n1794;
   wire n1795;
   wire n1796;
   wire n1797;
   wire n1798;
   wire n1799;
   wire n1800;
   wire n1801;
   wire n1802;
   wire n1803;
   wire n1804;
   wire n1805;
   wire n1806;
   wire n1807;
   wire n1808;
   wire n1809;
   wire n1810;
   wire n1811;
   wire n1812;
   wire n1813;
   wire n1814;
   wire n1815;
   wire n1816;
   wire n1817;
   wire n1818;
   wire n1819;
   wire n1820;
   wire n1821;
   wire n1822;
   wire n1823;
   wire n1824;
   wire n1825;
   wire n1826;
   wire n1827;
   wire n1828;
   wire n1829;
   wire n1830;
   wire n1831;
   wire n1832;
   wire n1833;
   wire n1834;
   wire n1835;
   wire n1836;
   wire n1837;
   wire n1838;
   wire n1839;
   wire n1840;
   wire n1841;
   wire n1842;
   wire n1843;
   wire n1844;
   wire n1845;
   wire n1846;
   wire n1847;
   wire n1848;
   wire n1849;
   wire n1850;
   wire n1851;
   wire n1852;
   wire n1853;
   wire n1854;
   wire n1855;
   wire n1856;
   wire n1857;
   wire n1858;
   wire n1859;
   wire n1860;
   wire n1861;
   wire n1862;
   wire n1863;
   wire n1864;
   wire n1865;
   wire n1866;
   wire n1867;
   wire n1868;
   wire n1869;
   wire n1870;
   wire n1871;
   wire n1872;
   wire n1873;
   wire n1874;
   wire n1875;
   wire n1876;
   wire n1877;
   wire n1878;
   wire n1879;
   wire n1880;
   wire n1881;
   wire n1882;
   wire n1883;
   wire n1884;
   wire n1885;
   wire n1886;
   wire n1887;
   wire n1888;
   wire n1889;
   wire n1890;
   wire n1891;
   wire n1892;
   wire n1893;
   wire n1894;
   wire n1895;
   wire n1896;
   wire n1897;
   wire n1898;
   wire n1899;
   wire n1900;
   wire n1901;
   wire n1902;
   wire n1903;
   wire n1904;
   wire n1905;
   wire n1906;
   wire n1907;
   wire n1908;
   wire n1909;
   wire n1910;
   wire n1911;
   wire n1912;
   wire n1913;
   wire n1914;
   wire n1915;
   wire n1916;
   wire n1917;
   wire n1918;
   wire n1919;
   wire n1920;
   wire n1921;
   wire n1922;
   wire n1923;
   wire n1924;
   wire n1925;
   wire n1926;
   wire n1927;
   wire n1928;
   wire n1929;
   wire n1930;
   wire n1931;
   wire n1932;
   wire n1933;
   wire n1934;
   wire n1935;
   wire n1936;
   wire n1937;
   wire n1938;
   wire n1939;
   wire n1940;
   wire n1941;
   wire n1942;
   wire n1943;
   wire n1944;
   wire n1945;
   wire n1946;
   wire n1947;
   wire n1948;
   wire n1949;
   wire n1950;
   wire n1951;
   wire n1952;
   wire n1953;
   wire n1954;
   wire n1955;
   wire n1956;
   wire n1957;
   wire n1958;
   wire n1959;
   wire n1960;
   wire n1961;
   wire n1962;
   wire n1963;
   wire n1964;
   wire n1965;
   wire n1966;
   wire n1967;
   wire n1968;
   wire n1969;
   wire n1970;
   wire n1971;
   wire n1972;
   wire n1973;
   wire n1974;
   wire n1975;
   wire n1976;
   wire n1977;
   wire n1978;
   wire n1979;
   wire n1980;
   wire n1981;
   wire n1982;
   wire n1983;
   wire n1984;
   wire n1985;
   wire n1986;
   wire n1987;
   wire n1988;
   wire n1989;
   wire n1990;
   wire n1991;
   wire n1992;
   wire n1993;
   wire n1994;
   wire n1995;
   wire n1996;
   wire n1997;
   wire n1998;
   wire n1999;
   wire n2000;
   wire n2001;
   wire n2002;
   wire n2003;
   wire n2004;
   wire n2005;
   wire n2006;
   wire n2007;
   wire n2008;
   wire n2009;
   wire n2010;
   wire n2011;
   wire n2012;
   wire n2013;
   wire n2014;
   wire n2015;
   wire n2016;
   wire n2017;
   wire n2018;
   wire n2019;
   wire n2020;
   wire n2021;
   wire n2022;
   wire n2023;
   wire n2024;
   wire n2025;
   wire n2026;
   wire n2027;
   wire n2028;
   wire n2029;
   wire n2030;
   wire n2031;
   wire n2032;
   wire n2033;
   wire n2034;
   wire n2035;
   wire n2036;
   wire n2037;
   wire n2038;
   wire n2039;
   wire n2040;
   wire n2041;
   wire n2042;
   wire n2043;
   wire n2044;
   wire n2045;
   wire n2046;
   wire n2047;
   wire n2048;
   wire n2049;
   wire n2050;
   wire n2051;
   wire n2052;
   wire n2053;
   wire n2054;
   wire n2055;
   wire n2056;
   wire n2057;
   wire n2058;
   wire n2059;
   wire n2060;
   wire n2061;
   wire n2062;
   wire n2063;
   wire n2064;
   wire n2065;
   wire n2066;
   wire n2067;
   wire n2068;
   wire n2069;
   wire n2070;
   wire n2071;
   wire n2072;
   wire n2073;
   wire n2074;
   wire n2075;
   wire n2076;
   wire n2077;
   wire n2078;
   wire n2079;
   wire n2080;
   wire n2081;
   wire n2082;
   wire n2083;
   wire n2084;
   wire n2085;
   wire n2086;
   wire n2087;
   wire n2088;
   wire n2089;
   wire n2090;
   wire n2091;
   wire n2092;
   wire n2093;
   wire n2094;
   wire n2095;
   wire n2096;
   wire n2097;
   wire n2098;
   wire n2099;
   wire n2100;
   wire n2101;
   wire n2102;
   wire n2103;
   wire n2104;
   wire n2105;
   wire n2106;
   wire n2107;
   wire n2108;
   wire n2109;
   wire n2110;
   wire n2111;
   wire n2112;
   wire n2113;
   wire n2114;
   wire n2115;
   wire n2116;
   wire n2117;
   wire n2118;
   wire n2119;
   wire n2120;
   wire n2121;
   wire n2122;
   wire n2123;
   wire n2124;
   wire n2125;
   wire n2126;
   wire n2127;
   wire n2128;
   wire n2129;
   wire n2130;
   wire n2131;
   wire n2132;
   wire n2133;
   wire n2134;
   wire n2135;
   wire n2136;
   wire n2137;
   wire n2138;
   wire n2139;
   wire n2140;
   wire n2141;
   wire n2142;
   wire n2143;
   wire n2144;
   wire n2145;
   wire n2146;
   wire n2147;
   wire n2148;
   wire n2149;
   wire n2150;
   wire n2151;
   wire n2152;
   wire n2153;
   wire n2154;
   wire n2155;
   wire n2156;
   wire n2157;
   wire n2158;
   wire n2159;
   wire n2160;
   wire n2161;
   wire n2162;
   wire n2163;
   wire n2164;
   wire n2165;
   wire n2166;
   wire n2167;
   wire n2168;
   wire n2169;
   wire n2170;
   wire n2171;
   wire n2172;
   wire n2173;
   wire n2174;
   wire n2175;
   wire n2176;
   wire n2177;
   wire n2178;
   wire n2179;
   wire n2180;
   wire n2181;
   wire n2182;
   wire n2183;
   wire n2184;
   wire n2185;
   wire n2186;
   wire n2187;
   wire n2188;
   wire n2189;
   wire n2190;
   wire n2191;
   wire n2192;
   wire n2193;
   wire n2194;
   wire n2195;
   wire n2196;
   wire n2197;
   wire n2198;
   wire n2199;
   wire n2200;
   wire n2201;
   wire n2202;
   wire n2203;
   wire n2204;
   wire n2205;
   wire n2206;
   wire n2207;
   wire n2208;
   wire n2209;
   wire n2210;
   wire n2211;
   wire n2212;
   wire n2213;
   wire n2214;
   wire n2215;
   wire n2216;
   wire n2217;
   wire n2218;
   wire n2219;
   wire n2220;
   wire n2221;
   wire n2222;
   wire n2223;
   wire n2224;
   wire n2225;
   wire n2226;
   wire n2227;
   wire n2228;
   wire n2229;
   wire n2230;
   wire n2231;
   wire n2232;
   wire n2233;
   wire n2234;
   wire n2235;
   wire n2236;
   wire n2237;
   wire n2238;
   wire n2239;
   wire n2240;
   wire n2241;
   wire n2242;
   wire n2243;
   wire n2244;
   wire n2245;
   wire n2246;
   wire n2247;
   wire n2248;
   wire n2249;
   wire n2250;
   wire n2251;
   wire n2252;
   wire n2253;
   wire n2254;
   wire n2255;
   wire n2256;
   wire n2257;
   wire n2258;
   wire n2259;
   wire n2260;
   wire n2261;
   wire n2262;
   wire n2263;
   wire n2264;
   wire n2265;
   wire n2266;
   wire n2267;
   wire n2268;
   wire n2269;
   wire n2270;
   wire n2271;
   wire n2272;
   wire n2273;
   wire n2274;
   wire n2275;
   wire n2276;
   wire n2277;
   wire n2278;
   wire n2279;
   wire n2280;
   wire n2281;
   wire n2282;
   wire n2283;
   wire n2284;
   wire n2285;
   wire n2286;
   wire n2287;
   wire n2288;
   wire n2289;
   wire n2290;
   wire n2291;
   wire n2292;
   wire n2293;
   wire n2294;
   wire n2295;
   wire n2296;
   wire n2297;
   wire n2298;
   wire n2299;
   wire n2300;
   wire n2301;
   wire n2302;
   wire n2303;
   wire n2304;
   wire n2305;
   wire n2306;
   wire n2307;
   wire n2308;
   wire n2309;
   wire n2310;
   wire n2311;
   wire n2312;
   wire n2313;
   wire n2314;
   wire n2315;
   wire n2316;
   wire n2317;
   wire n2318;
   wire n2319;
   wire n2320;
   wire n2321;
   wire n2322;
   wire n2323;
   wire n2324;
   wire n2325;
   wire n2326;
   wire n2327;
   wire n2328;
   wire n2329;
   wire n2330;
   wire n2331;
   wire n2332;
   wire n2333;
   wire n2334;
   wire n2335;
   wire n2336;
   wire n2337;
   wire n2338;
   wire n2339;
   wire n2340;
   wire n2341;
   wire n2342;
   wire n2343;
   wire n2344;
   wire n2345;
   wire n2346;
   wire n2347;
   wire n2348;
   wire n2349;
   wire n2350;
   wire n2351;
   wire n2352;
   wire n2353;
   wire n2354;
   wire n2355;
   wire n2356;
   wire n2357;
   wire n2358;
   wire n2359;
   wire n2360;
   wire n2361;
   wire n2362;
   wire n2363;
   wire n2364;
   wire n2365;
   wire n2366;
   wire n2367;
   wire n2368;
   wire n2369;
   wire n2370;
   wire n2371;
   wire n2372;
   wire n2373;
   wire n2374;
   wire n2375;
   wire n2376;
   wire n2377;
   wire n2378;
   wire n2379;
   wire n2380;
   wire n2381;
   wire n2382;
   wire n2383;
   wire n2384;
   wire n2385;
   wire n2386;
   wire n2387;
   wire n2388;
   wire n2389;
   wire n2390;
   wire n2391;
   wire n2392;
   wire n2393;
   wire n2394;
   wire n2395;
   wire n2396;
   wire n2397;
   wire n2398;
   wire n2399;
   wire n2400;
   wire n2401;
   wire n2402;
   wire n2403;
   wire n2404;
   wire n2405;
   wire n2406;
   wire n2407;
   wire n2408;
   wire n2409;
   wire n2410;
   wire n2411;
   wire n2412;
   wire n2413;
   wire n2414;
   wire n2415;
   wire n2416;
   wire n2417;
   wire n2418;
   wire n2419;
   wire n2420;
   wire n2421;
   wire n2422;
   wire n2423;
   wire n2424;
   wire n2425;
   wire n2426;
   wire n2427;
   wire n2428;
   wire n2429;
   wire n2430;
   wire n2431;
   wire n2432;
   wire n2433;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n7;
   wire n8;
   wire n2622;
   wire n2623;
   wire n2624;
   wire n2637;
   wire n2638;
   wire n2639;
   wire n2640;
   wire n2641;
   wire n2642;
   wire n2643;
   wire n2644;
   wire n2645;
   wire n2646;
   wire n2647;
   wire n2648;
   wire n2649;
   wire n2650;
   wire n2651;
   wire n2652;
   wire n2653;
   wire n2654;
   wire n2655;
   wire n2656;
   wire n2657;
   wire n2658;
   wire n2659;
   wire n2660;
   wire n2661;
   wire n2662;
   wire n2663;
   wire n2664;
   wire n2665;
   wire n2666;
   wire n2667;
   wire n2668;
   wire n2669;
   wire n2670;
   wire n2671;
   wire n2672;
   wire n2673;
   wire n2674;
   wire n2675;
   wire n2676;
   wire n2677;
   wire n2678;
   wire n2679;
   wire n2680;
   wire n2681;
   wire n2682;
   wire n2683;
   wire n2684;
   wire n2685;
   wire n2686;
   wire n2687;
   wire n2688;
   wire n2689;
   wire n2690;
   wire n2691;
   wire n2692;
   wire n2693;
   wire n2694;
   wire n2695;
   wire n2696;
   wire n2697;
   wire n2698;
   wire n2699;
   wire n2766;
   wire n2769;
   wire n2770;
   wire n2773;
   wire n2775;
   wire n2780;
   wire n2781;
   wire n2784;
   wire n2800;
   wire n2806;
   wire n2817;
   wire n2818;
   wire n2823;
   wire n2824;
   wire n2827;
   wire n2828;
   wire n2829;
   wire n2868;
   wire n2869;
   wire n2870;
   wire n2871;
   wire n2872;
   wire n2873;
   wire n2874;
   wire n2875;
   wire n2876;
   wire n2877;
   wire n2878;
   wire n2879;
   wire [1407:0] key_mem;
   wire [7:0] rcon_reg;
   wire [1:0] key_mem_ctrl_reg;
   wire [3:0] round_ctr_reg;
   wire [127:32] prev_key1_reg;

   BUFXL FE_PHC5077_n2415 (.Y(FE_PHN5077_n2415), 
	.A(FE_PHN5065_n2415));
   BUFXL FE_PHC5076_n2407 (.Y(FE_PHN5076_n2407), 
	.A(FE_PHN5066_n2407));
   CLKBUFX1 FE_PHC5073_n2430 (.Y(FE_PHN5073_n2430), 
	.A(FE_PHN3409_n2430));
   CLKBUFX1 FE_PHC5066_n2407 (.Y(FE_PHN5066_n2407), 
	.A(n2407));
   CLKBUFX3 FE_PHC5065_n2415 (.Y(FE_PHN5065_n2415), 
	.A(n2415));
   DLY2X1 FE_PHC5063_n2400 (.Y(FE_PHN5063_n2400), 
	.A(n2400));
   DLY2X1 FE_PHC5062_n2416 (.Y(FE_PHN5062_n2416), 
	.A(n2416));
   DLY2X1 FE_PHC5061_n2391 (.Y(FE_PHN5061_n2391), 
	.A(n2391));
   DLY2X1 FE_PHC5060_n2408 (.Y(FE_PHN5060_n2408), 
	.A(n2408));
   DLY2X1 FE_PHC5058_n2392 (.Y(FE_PHN5058_n2392), 
	.A(n2392));
   DLY2X1 FE_PHC5057_n2399 (.Y(FE_PHN5057_n2399), 
	.A(n2399));
   DLY2X1 FE_PHC5056_n2412 (.Y(FE_PHN5056_n2412), 
	.A(n2412));
   DLY2X1 FE_PHC5055_n2409 (.Y(FE_PHN5055_n2409), 
	.A(n2409));
   DLY2X1 FE_PHC5054_n2403 (.Y(FE_PHN5054_n2403), 
	.A(n2403));
   DLY2X1 FE_PHC5053_n2393 (.Y(FE_PHN5053_n2393), 
	.A(n2393));
   DLY2X1 FE_PHC5052_n2417 (.Y(FE_PHN5052_n2417), 
	.A(n2417));
   DLY2X1 FE_PHC5051_n2404 (.Y(FE_PHN5051_n2404), 
	.A(n2404));
   DLY2X1 FE_PHC5050_n2411 (.Y(FE_PHN5050_n2411), 
	.A(n2411));
   DLY2X1 FE_PHC5049_n2401 (.Y(FE_PHN5049_n2401), 
	.A(n2401));
   DLY2X1 FE_PHC5047_n2431 (.Y(FE_PHN5047_n2431), 
	.A(n2431));
   DLY2X1 FE_PHC5044_n2397 (.Y(FE_PHN5044_n2397), 
	.A(n2397));
   DLY2X1 FE_PHC5043_n2406 (.Y(FE_PHN5043_n2406), 
	.A(n2406));
   DLY2X1 FE_PHC5042_n2394 (.Y(FE_PHN5042_n2394), 
	.A(n2394));
   DLY2X1 FE_PHC5041_n2398 (.Y(FE_PHN5041_n2398), 
	.A(n2398));
   DLY2X1 FE_PHC5040_n2410 (.Y(FE_PHN5040_n2410), 
	.A(n2410));
   DLY2X1 FE_PHC5039_n2405 (.Y(FE_PHN5039_n2405), 
	.A(n2405));
   DLY4X1 FE_PHC5038_n2420 (.Y(FE_PHN5038_n2420), 
	.A(n2420));
   DLY2X1 FE_PHC5037_n2402 (.Y(FE_PHN5037_n2402), 
	.A(n2402));
   DLY4X1 FE_PHC5036_n2359 (.Y(FE_PHN5036_n2359), 
	.A(n2359));
   DLY4X1 FE_PHC5035_n2419 (.Y(FE_PHN5035_n2419), 
	.A(n2419));
   DLY4X1 FE_PHC5034_n2351 (.Y(FE_PHN5034_n2351), 
	.A(n2351));
   DLY3X1 FE_PHC5033_n2414 (.Y(FE_PHN5033_n2414), 
	.A(n2414));
   DLY4X1 FE_PHC5032_n2390 (.Y(FE_PHN5032_n2390), 
	.A(n2390));
   DLY3X1 FE_PHC5031_n2413 (.Y(FE_PHN5031_n2413), 
	.A(n2413));
   DLY4X1 FE_PHC5030_n2418 (.Y(FE_PHN5030_n2418), 
	.A(n2418));
   DLY3X1 FE_PHC5029_n2352 (.Y(FE_PHN5029_n2352), 
	.A(n2352));
   DLY4X1 FE_PHC5028_n2363 (.Y(FE_PHN5028_n2363), 
	.A(n2363));
   DLY3X1 FE_PHC5027_n2396 (.Y(FE_PHN5027_n2396), 
	.A(n2396));
   DLY3X1 FE_PHC5026_n2353 (.Y(FE_PHN5026_n2353), 
	.A(n2353));
   DLY3X1 FE_PHC5025_n2354 (.Y(FE_PHN5025_n2354), 
	.A(n2354));
   DLY3X1 FE_PHC5024_n2344 (.Y(FE_PHN5024_n2344), 
	.A(n2344));
   DLY4X1 FE_PHC5023_n2293 (.Y(FE_PHN5023_n2293), 
	.A(n2293));
   DLY3X1 FE_PHC5022_n2356 (.Y(FE_PHN5022_n2356), 
	.A(n2356));
   DLY3X1 FE_PHC5021_n2297 (.Y(FE_PHN5021_n2297), 
	.A(n2297));
   DLY4X1 FE_PHC5020_n2395 (.Y(FE_PHN5020_n2395), 
	.A(n2395));
   DLY4X1 FE_PHC5019_n2349 (.Y(FE_PHN5019_n2349), 
	.A(n2349));
   DLY3X1 FE_PHC5018_n2300 (.Y(FE_PHN5018_n2300), 
	.A(n2300));
   DLY3X1 FE_PHC5017_n2362 (.Y(FE_PHN5017_n2362), 
	.A(n2362));
   DLY3X1 FE_PHC5016_n2335 (.Y(FE_PHN5016_n2335), 
	.A(n2335));
   DLY4X1 FE_PHC5015_n2360 (.Y(FE_PHN5015_n2360), 
	.A(n2360));
   DLY4X1 FE_PHC5014_n2295 (.Y(FE_PHN5014_n2295), 
	.A(n2295));
   DLY4X1 FE_PHC5013_n2346 (.Y(FE_PHN5013_n2346), 
	.A(n2346));
   DLY4X1 FE_PHC5012_n2345 (.Y(FE_PHN5012_n2345), 
	.A(n2345));
   DLY3X1 FE_PHC5011_n2336 (.Y(FE_PHN5011_n2336), 
	.A(n2336));
   DLY3X1 FE_PHC5010_n2357 (.Y(FE_PHN5010_n2357), 
	.A(n2357));
   DLY3X1 FE_PHC5009_n2361 (.Y(FE_PHN5009_n2361), 
	.A(n2361));
   DLY4X1 FE_PHC5008_n2348 (.Y(FE_PHN5008_n2348), 
	.A(n2348));
   DLY4X1 FE_PHC5007_n2341 (.Y(FE_PHN5007_n2341), 
	.A(n2341));
   DLY4X1 FE_PHC5006_n2364 (.Y(FE_PHN5006_n2364), 
	.A(n2364));
   DLY3X1 FE_PHC5005_n2296 (.Y(FE_PHN5005_n2296), 
	.A(n2296));
   DLY3X1 FE_PHC5004_n2339 (.Y(FE_PHN5004_n2339), 
	.A(n2339));
   DLY3X1 FE_PHC5003_n2340 (.Y(FE_PHN5003_n2340), 
	.A(n2340));
   DLY3X1 FE_PHC5002_n2347 (.Y(FE_PHN5002_n2347), 
	.A(n2347));
   DLY4X1 FE_PHC5001_n2342 (.Y(FE_PHN5001_n2342), 
	.A(n2342));
   DLY4X1 FE_PHC5000_n2343 (.Y(FE_PHN5000_n2343), 
	.A(n2343));
   DLY4X1 FE_PHC4999_n2338 (.Y(FE_PHN4999_n2338), 
	.A(n2338));
   DLY4X1 FE_PHC4998_n2355 (.Y(FE_PHN4998_n2355), 
	.A(n2355));
   DLY3X1 FE_PHC4997_n2389 (.Y(FE_PHN4997_n2389), 
	.A(n2389));
   DLY3X1 FE_PHC4996_key_mem_846_ (.Y(FE_PHN4996_key_mem_846_), 
	.A(key_mem[846]));
   DLY4X1 FE_PHC4995_n2334 (.Y(FE_PHN4995_n2334), 
	.A(n2334));
   DLY3X1 FE_PHC4994_n2358 (.Y(FE_PHN4994_n2358), 
	.A(n2358));
   DLY3X1 FE_PHC4993_n2294 (.Y(FE_PHN4993_n2294), 
	.A(n2294));
   DLY3X1 FE_PHC4992_n2299 (.Y(FE_PHN4992_n2299), 
	.A(n2299));
   DLY4X1 FE_PHC4991_n1210 (.Y(FE_PHN4991_n1210), 
	.A(n1210));
   DLY3X1 FE_PHC4990_n2333 (.Y(FE_PHN4990_n2333), 
	.A(n2333));
   DLY3X1 FE_PHC4989_n2337 (.Y(FE_PHN4989_n2337), 
	.A(n2337));
   DLY4X1 FE_PHC4988_n1730 (.Y(FE_PHN4988_n1730), 
	.A(n1730));
   DLY4X1 FE_PHC4987_n1916 (.Y(FE_PHN4987_n1916), 
	.A(n1916));
   DLY4X1 FE_PHC4986_n2298 (.Y(FE_PHN4986_n2298), 
	.A(n2298));
   DLY3X1 FE_PHC4985_n1981 (.Y(FE_PHN4985_n1981), 
	.A(n1981));
   DLY3X1 FE_PHC4984_n2350 (.Y(FE_PHN4984_n2350), 
	.A(n2350));
   DLY3X1 FE_PHC4983_n1052 (.Y(FE_PHN4983_n1052), 
	.A(n1052));
   DLY3X1 FE_PHC4982_n1207 (.Y(FE_PHN4982_n1207), 
	.A(n1207));
   DLY3X1 FE_PHC4981_n1178 (.Y(FE_PHN4981_n1178), 
	.A(n1178));
   DLY3X1 FE_PHC4980_n2425 (.Y(FE_PHN4980_n2425), 
	.A(n2425));
   DLY4X1 FE_PHC4979_n1085 (.Y(FE_PHN4979_n1085), 
	.A(n1085));
   DLY4X1 FE_PHC4978_n1027 (.Y(FE_PHN4978_n1027), 
	.A(n1027));
   DLY4X1 FE_PHC4977_n1329 (.Y(FE_PHN4977_n1329), 
	.A(n1329));
   DLY4X1 FE_PHC4976_n1239 (.Y(FE_PHN4976_n1239), 
	.A(n1239));
   DLY3X1 FE_PHC4975_n1246 (.Y(FE_PHN4975_n1246), 
	.A(n1246));
   DLY4X1 FE_PHC4974_n1192 (.Y(FE_PHN4974_n1192), 
	.A(n1192));
   DLY4X1 FE_PHC4973_n2304 (.Y(FE_PHN4973_n2304), 
	.A(n2304));
   DLY4X1 FE_PHC4972_n1224 (.Y(FE_PHN4972_n1224), 
	.A(n1224));
   DLY4X1 FE_PHC4971_n1020 (.Y(FE_PHN4971_n1020), 
	.A(n1020));
   DLY3X1 FE_PHC4970_n957 (.Y(FE_PHN4970_n957), 
	.A(n957));
   DLY4X1 FE_PHC4969_n1116 (.Y(FE_PHN4969_n1116), 
	.A(n1116));
   DLY4X1 FE_PHC4968_n2312 (.Y(FE_PHN4968_n2312), 
	.A(n2312));
   DLY4X1 FE_PHC4967_n1179 (.Y(FE_PHN4967_n1179), 
	.A(n1179));
   DLY4X1 FE_PHC4966_n1067 (.Y(FE_PHN4966_n1067), 
	.A(n1067));
   DLY4X1 FE_PHC4965_n918 (.Y(FE_PHN4965_n918), 
	.A(n918));
   DLY3X1 FE_PHC4964_n1558 (.Y(FE_PHN4964_n1558), 
	.A(n1558));
   DLY3X1 FE_PHC4963_n1073 (.Y(FE_PHN4963_n1073), 
	.A(n1073));
   DLY3X1 FE_PHC4961_n1191 (.Y(FE_PHN4961_n1191), 
	.A(n1191));
   DLY3X1 FE_PHC4960_n1118 (.Y(FE_PHN4960_n1118), 
	.A(n1118));
   DLY4X1 FE_PHC4959_n1033 (.Y(FE_PHN4959_n1033), 
	.A(n1033));
   DLY4X1 FE_PHC4958_n1062 (.Y(FE_PHN4958_n1062), 
	.A(n1062));
   DLY4X1 FE_PHC4956_n1319 (.Y(FE_PHN4956_n1319), 
	.A(n1319));
   DLY4X1 FE_PHC4955_n1390 (.Y(FE_PHN4955_n1390), 
	.A(n1390));
   DLY3X1 FE_PHC4954_n2376 (.Y(FE_PHN4954_n2376), 
	.A(n2376));
   DLY3X1 FE_PHC4953_n1978 (.Y(FE_PHN4953_n1978), 
	.A(n1978));
   DLY3X1 FE_PHC4952_n931 (.Y(FE_PHN4952_n931), 
	.A(n931));
   DLY3X1 FE_PHC4951_n1263 (.Y(FE_PHN4951_n1263), 
	.A(n1263));
   DLY4X1 FE_PHC4950_n1612 (.Y(FE_PHN4950_n1612), 
	.A(n1612));
   DLY4X1 FE_PHC4949_n1231 (.Y(FE_PHN4949_n1231), 
	.A(n1231));
   DLY4X1 FE_PHC4948_n2379 (.Y(FE_PHN4948_n2379), 
	.A(n2379));
   DLY3X1 FE_PHC4947_n1359 (.Y(FE_PHN4947_n1359), 
	.A(n1359));
   DLY3X1 FE_PHC4946_n1208 (.Y(FE_PHN4946_n1208), 
	.A(n1208));
   DLY3X1 FE_PHC4945_n1327 (.Y(FE_PHN4945_n1327), 
	.A(n1327));
   DLY3X1 FE_PHC4944_n1268 (.Y(FE_PHN4944_n1268), 
	.A(n1268));
   DLY3X1 FE_PHC4943_n1243 (.Y(FE_PHN4943_n1243), 
	.A(n1243));
   DLY3X1 FE_PHC4942_n2385 (.Y(FE_PHN4942_n2385), 
	.A(n2385));
   DLY4X1 FE_PHC4941_n1932 (.Y(FE_PHN4941_n1932), 
	.A(n1932));
   DLY4X1 FE_PHC4940_n2370 (.Y(FE_PHN4940_n2370), 
	.A(n2370));
   DLY4X1 FE_PHC4939_n965 (.Y(FE_PHN4939_n965), 
	.A(n965));
   DLY4X1 FE_PHC4938_n992 (.Y(FE_PHN4938_n992), 
	.A(n992));
   DLY4X1 FE_PHC4937_n1248 (.Y(FE_PHN4937_n1248), 
	.A(n1248));
   DLY4X1 FE_PHC4936_n1308 (.Y(FE_PHN4936_n1308), 
	.A(n1308));
   DLY4X1 FE_PHC4935_n1099 (.Y(FE_PHN4935_n1099), 
	.A(n1099));
   DLY4X1 FE_PHC4934_n1173 (.Y(FE_PHN4934_n1173), 
	.A(n1173));
   DLY4X1 FE_PHC4933_n1537 (.Y(FE_PHN4933_n1537), 
	.A(n1537));
   DLY3X1 FE_PHC4932_n1126 (.Y(FE_PHN4932_n1126), 
	.A(n1126));
   DLY3X1 FE_PHC4931_n981 (.Y(FE_PHN4931_n981), 
	.A(n981));
   DLY3X1 FE_PHC4930_n1571 (.Y(FE_PHN4930_n1571), 
	.A(n1571));
   DLY4X1 FE_PHC4929_n1233 (.Y(FE_PHN4929_n1233), 
	.A(n1233));
   DLY3X1 FE_PHC4928_n2091 (.Y(FE_PHN4928_n2091), 
	.A(FE_PHN2755_n2091));
   DLY3X1 FE_PHC4927_n1621 (.Y(FE_PHN4927_n1621), 
	.A(n1621));
   DLY3X1 FE_PHC4926_n1261 (.Y(FE_PHN4926_n1261), 
	.A(n1261));
   DLY3X1 FE_PHC4925_n1038 (.Y(FE_PHN4925_n1038), 
	.A(n1038));
   DLY3X1 FE_PHC4924_n1209 (.Y(FE_PHN4924_n1209), 
	.A(n1209));
   DLY4X1 FE_PHC4923_n1154 (.Y(FE_PHN4923_n1154), 
	.A(n1154));
   DLY4X1 FE_PHC4922_n1252 (.Y(FE_PHN4922_n1252), 
	.A(n1252));
   DLY4X1 FE_PHC4921_n1267 (.Y(FE_PHN4921_n1267), 
	.A(n1267));
   DLY4X1 FE_PHC4920_n1599 (.Y(FE_PHN4920_n1599), 
	.A(n1599));
   DLY4X1 FE_PHC4919_n1152 (.Y(FE_PHN4919_n1152), 
	.A(n1152));
   DLY4X1 FE_PHC4918_n1999 (.Y(FE_PHN4918_n1999), 
	.A(n1999));
   DLY4X1 FE_PHC4917_n1247 (.Y(FE_PHN4917_n1247), 
	.A(n1247));
   DLY4X1 FE_PHC4916_n1193 (.Y(FE_PHN4916_n1193), 
	.A(n1193));
   DLY3X1 FE_PHC4915_n1180 (.Y(FE_PHN4915_n1180), 
	.A(n1180));
   DLY4X1 FE_PHC4914_n1933 (.Y(FE_PHN4914_n1933), 
	.A(n1933));
   DLY3X1 FE_PHC4913_n1048 (.Y(FE_PHN4913_n1048), 
	.A(n1048));
   DLY3X1 FE_PHC4912_n1262 (.Y(FE_PHN4912_n1262), 
	.A(n1262));
   DLY3X1 FE_PHC4911_n1253 (.Y(FE_PHN4911_n1253), 
	.A(n1253));
   DLY3X1 FE_PHC4910_n1888 (.Y(FE_PHN4910_n1888), 
	.A(n1888));
   DLY3X1 FE_PHC4909_n1149 (.Y(FE_PHN4909_n1149), 
	.A(n1149));
   DLY4X1 FE_PHC4908_n1141 (.Y(FE_PHN4908_n1141), 
	.A(n1141));
   DLY4X1 FE_PHC4907_n1256 (.Y(FE_PHN4907_n1256), 
	.A(n1256));
   DLY3X1 FE_PHC4906_n1142 (.Y(FE_PHN4906_n1142), 
	.A(n1142));
   DLY3X1 FE_PHC4905_n1607 (.Y(FE_PHN4905_n1607), 
	.A(n1607));
   DLY3X1 FE_PHC4904_n1137 (.Y(FE_PHN4904_n1137), 
	.A(n1137));
   DLY3X1 FE_PHC4903_n1194 (.Y(FE_PHN4903_n1194), 
	.A(n1194));
   DLY4X1 FE_PHC4902_n1214 (.Y(FE_PHN4902_n1214), 
	.A(n1214));
   DLY4X1 FE_PHC4901_n1886 (.Y(FE_PHN4901_n1886), 
	.A(n1886));
   DLY4X1 FE_PHC4900_n1220 (.Y(FE_PHN4900_n1220), 
	.A(n1220));
   DLY4X1 FE_PHC4899_n2365 (.Y(FE_PHN4899_n2365), 
	.A(n2365));
   DLY4X1 FE_PHC4898_n1037 (.Y(FE_PHN4898_n1037), 
	.A(n1037));
   DLY4X1 FE_PHC4897_n974 (.Y(FE_PHN4897_n974), 
	.A(n974));
   DLY4X1 FE_PHC4896_n958 (.Y(FE_PHN4896_n958), 
	.A(n958));
   DLY4X1 FE_PHC4895_n2428 (.Y(FE_PHN4895_n2428), 
	.A(n2428));
   DLY4X1 FE_PHC4894_n1984 (.Y(FE_PHN4894_n1984), 
	.A(n1984));
   DLY4X1 FE_PHC4893_n1186 (.Y(FE_PHN4893_n1186), 
	.A(n1186));
   DLY4X1 FE_PHC4892_n1221 (.Y(FE_PHN4892_n1221), 
	.A(n1221));
   DLY4X1 FE_PHC4891_n1198 (.Y(FE_PHN4891_n1198), 
	.A(n1198));
   DLY4X1 FE_PHC4890_n1139 (.Y(FE_PHN4890_n1139), 
	.A(n1139));
   DLY4X1 FE_PHC4889_n1086 (.Y(FE_PHN4889_n1086), 
	.A(n1086));
   DLY4X1 FE_PHC4888_n2327 (.Y(FE_PHN4888_n2327), 
	.A(n2327));
   DLY4X1 FE_PHC4887_n1371 (.Y(FE_PHN4887_n1371), 
	.A(n1371));
   DLY4X1 FE_PHC4886_n1293 (.Y(FE_PHN4886_n1293), 
	.A(n1293));
   DLY3X1 FE_PHC4885_n2229 (.Y(FE_PHN4885_n2229), 
	.A(n2229));
   DLY3X1 FE_PHC4884_n2313 (.Y(FE_PHN4884_n2313), 
	.A(n2313));
   DLY4X1 FE_PHC4883_n2017 (.Y(FE_PHN4883_n2017), 
	.A(n2017));
   DLY3X1 FE_PHC4882_n1144 (.Y(FE_PHN4882_n1144), 
	.A(n1144));
   DLY3X1 FE_PHC4881_n1586 (.Y(FE_PHN4881_n1586), 
	.A(n1586));
   DLY3X1 FE_PHC4880_n1001 (.Y(FE_PHN4880_n1001), 
	.A(n1001));
   DLY3X1 FE_PHC4879_n1232 (.Y(FE_PHN4879_n1232), 
	.A(n1232));
   DLY3X1 FE_PHC4878_n1244 (.Y(FE_PHN4878_n1244), 
	.A(n1244));
   DLY3X1 FE_PHC4877_n1965 (.Y(FE_PHN4877_n1965), 
	.A(n1965));
   DLY3X1 FE_PHC4876_n2319 (.Y(FE_PHN4876_n2319), 
	.A(n2319));
   DLY3X1 FE_PHC4875_n1989 (.Y(FE_PHN4875_n1989), 
	.A(n1989));
   DLY3X1 FE_PHC4874_n2326 (.Y(FE_PHN4874_n2326), 
	.A(n2326));
   DLY3X1 FE_PHC4873_n1021 (.Y(FE_PHN4873_n1021), 
	.A(n1021));
   DLY4X1 FE_PHC4872_n1344 (.Y(FE_PHN4872_n1344), 
	.A(n1344));
   DLY4X1 FE_PHC4871_n886 (.Y(FE_PHN4871_n886), 
	.A(n886));
   DLY4X1 FE_PHC4870_n1045 (.Y(FE_PHN4870_n1045), 
	.A(n1045));
   DLY4X1 FE_PHC4869_n1976 (.Y(FE_PHN4869_n1976), 
	.A(n1976));
   DLY4X1 FE_PHC4868_n1563 (.Y(FE_PHN4868_n1563), 
	.A(n1563));
   DLY4X1 FE_PHC4867_n1393 (.Y(FE_PHN4867_n1393), 
	.A(n1393));
   DLY4X1 FE_PHC4866_n1943 (.Y(FE_PHN4866_n1943), 
	.A(n1943));
   DLY4X1 FE_PHC4865_n1356 (.Y(FE_PHN4865_n1356), 
	.A(n1356));
   DLY4X1 FE_PHC4864_n1598 (.Y(FE_PHN4864_n1598), 
	.A(n1598));
   DLY4X1 FE_PHC4863_n1526 (.Y(FE_PHN4863_n1526), 
	.A(n1526));
   DLY4X1 FE_PHC4862_n1106 (.Y(FE_PHN4862_n1106), 
	.A(n1106));
   DLY4X1 FE_PHC4861_n1827 (.Y(FE_PHN4861_n1827), 
	.A(n1827));
   DLY4X1 FE_PHC4860_n1087 (.Y(FE_PHN4860_n1087), 
	.A(n1087));
   DLY4X1 FE_PHC4859_n935 (.Y(FE_PHN4859_n935), 
	.A(n935));
   DLY4X1 FE_PHC4858_n1264 (.Y(FE_PHN4858_n1264), 
	.A(n1264));
   DLY3X1 FE_PHC4857_n1304 (.Y(FE_PHN4857_n1304), 
	.A(n1304));
   DLY3X1 FE_PHC4856_n1189 (.Y(FE_PHN4856_n1189), 
	.A(n1189));
   DLY4X1 FE_PHC4855_n1230 (.Y(FE_PHN4855_n1230), 
	.A(n1230));
   DLY4X1 FE_PHC4853_n1158 (.Y(FE_PHN4853_n1158), 
	.A(n1158));
   DLY4X1 FE_PHC4852_n1649 (.Y(FE_PHN4852_n1649), 
	.A(n1649));
   DLY3X1 FE_PHC4851_n2371 (.Y(FE_PHN4851_n2371), 
	.A(n2371));
   DLY3X1 FE_PHC4850_n1203 (.Y(FE_PHN4850_n1203), 
	.A(n1203));
   DLY3X1 FE_PHC4849_n2035 (.Y(FE_PHN4849_n2035), 
	.A(n2035));
   DLY3X1 FE_PHC4848_n1165 (.Y(FE_PHN4848_n1165), 
	.A(n1165));
   DLY3X1 FE_PHC4847_n1009 (.Y(FE_PHN4847_n1009), 
	.A(n1009));
   DLY4X1 FE_PHC4846_n1115 (.Y(FE_PHN4846_n1115), 
	.A(n1115));
   DLY3X1 FE_PHC4845_n2315 (.Y(FE_PHN4845_n2315), 
	.A(n2315));
   DLY3X1 FE_PHC4844_n1647 (.Y(FE_PHN4844_n1647), 
	.A(n1647));
   DLY3X1 FE_PHC4843_n1228 (.Y(FE_PHN4843_n1228), 
	.A(n1228));
   DLY4X1 FE_PHC4842_n1251 (.Y(FE_PHN4842_n1251), 
	.A(n1251));
   DLY3X1 FE_PHC4841_n1134 (.Y(FE_PHN4841_n1134), 
	.A(n1134));
   DLY4X1 FE_PHC4840_n2332 (.Y(FE_PHN4840_n2332), 
	.A(n2332));
   DLY4X1 FE_PHC4839_n1872 (.Y(FE_PHN4839_n1872), 
	.A(n1872));
   DLY4X1 FE_PHC4838_n1282 (.Y(FE_PHN4838_n1282), 
	.A(n1282));
   DLY4X1 FE_PHC4837_n1171 (.Y(FE_PHN4837_n1171), 
	.A(n1171));
   DLY4X1 FE_PHC4836_n1501 (.Y(FE_PHN4836_n1501), 
	.A(FE_PHN2727_n1501));
   DLY4X1 FE_PHC4835_n2036 (.Y(FE_PHN4835_n2036), 
	.A(n2036));
   DLY4X1 FE_PHC4834_n1070 (.Y(FE_PHN4834_n1070), 
	.A(n1070));
   DLY4X1 FE_PHC4833_n1630 (.Y(FE_PHN4833_n1630), 
	.A(n1630));
   DLY4X1 FE_PHC4832_n1617 (.Y(FE_PHN4832_n1617), 
	.A(n1617));
   DLY4X1 FE_PHC4831_n1100 (.Y(FE_PHN4831_n1100), 
	.A(n1100));
   DLY4X1 FE_PHC4830_n1614 (.Y(FE_PHN4830_n1614), 
	.A(n1614));
   DLY4X1 FE_PHC4829_n1223 (.Y(FE_PHN4829_n1223), 
	.A(n1223));
   DLY4X1 FE_PHC4828_n1608 (.Y(FE_PHN4828_n1608), 
	.A(n1608));
   DLY4X1 FE_PHC4827_n954 (.Y(FE_PHN4827_n954), 
	.A(n954));
   DLY4X1 FE_PHC4826_n1065 (.Y(FE_PHN4826_n1065), 
	.A(n1065));
   DLY4X1 FE_PHC4825_n1632 (.Y(FE_PHN4825_n1632), 
	.A(n1632));
   DLY4X1 FE_PHC4824_n1172 (.Y(FE_PHN4824_n1172), 
	.A(n1172));
   DLY4X1 FE_PHC4823_n1204 (.Y(FE_PHN4823_n1204), 
	.A(n1204));
   DLY4X1 FE_PHC4822_n1091 (.Y(FE_PHN4822_n1091), 
	.A(n1091));
   DLY3X1 FE_PHC4821_n1962 (.Y(FE_PHN4821_n1962), 
	.A(n1962));
   DLY3X1 FE_PHC4820_n1199 (.Y(FE_PHN4820_n1199), 
	.A(n1199));
   DLY3X1 FE_PHC4819_n1148 (.Y(FE_PHN4819_n1148), 
	.A(n1148));
   DLY3X1 FE_PHC4818_n1973 (.Y(FE_PHN4818_n1973), 
	.A(n1973));
   DLY3X1 FE_PHC4817_n1348 (.Y(FE_PHN4817_n1348), 
	.A(n1348));
   DLY3X1 FE_PHC4816_n1249 (.Y(FE_PHN4816_n1249), 
	.A(n1249));
   DLY4X1 FE_PHC4815_n1156 (.Y(FE_PHN4815_n1156), 
	.A(n1156));
   DLY3X1 FE_PHC4814_n2308 (.Y(FE_PHN4814_n2308), 
	.A(n2308));
   DLY3X1 FE_PHC4813_n1355 (.Y(FE_PHN4813_n1355), 
	.A(n1355));
   DLY3X1 FE_PHC4812_n2302 (.Y(FE_PHN4812_n2302), 
	.A(n2302));
   DLY3X1 FE_PHC4811_n1241 (.Y(FE_PHN4811_n1241), 
	.A(n1241));
   DLY4X1 FE_PHC4810_n1557 (.Y(FE_PHN4810_n1557), 
	.A(n1557));
   DLY3X1 FE_PHC4809_n2366 (.Y(FE_PHN4809_n2366), 
	.A(n2366));
   DLY3X1 FE_PHC4808_n1488 (.Y(FE_PHN4808_n1488), 
	.A(n1488));
   DLY3X1 FE_PHC4807_n1681 (.Y(FE_PHN4807_n1681), 
	.A(n1681));
   DLY4X1 FE_PHC4806_n1619 (.Y(FE_PHN4806_n1619), 
	.A(n1619));
   DLY3X1 FE_PHC4805_n1300 (.Y(FE_PHN4805_n1300), 
	.A(n1300));
   DLY4X1 FE_PHC4804_n1039 (.Y(FE_PHN4804_n1039), 
	.A(n1039));
   DLY4X1 FE_PHC4803_n1587 (.Y(FE_PHN4803_n1587), 
	.A(n1587));
   DLY3X1 FE_PHC4802_n1611 (.Y(FE_PHN4802_n1611), 
	.A(n1611));
   DLY3X1 FE_PHC4801_n1307 (.Y(FE_PHN4801_n1307), 
	.A(n1307));
   DLY3X1 FE_PHC4800_n1066 (.Y(FE_PHN4800_n1066), 
	.A(n1066));
   DLY3X1 FE_PHC4799_n1326 (.Y(FE_PHN4799_n1326), 
	.A(n1326));
   DLY3X1 FE_PHC4798_n969 (.Y(FE_PHN4798_n969), 
	.A(n969));
   DLY4X1 FE_PHC4797_n1561 (.Y(FE_PHN4797_n1561), 
	.A(n1561));
   DLY3X1 FE_PHC4796_n1206 (.Y(FE_PHN4796_n1206), 
	.A(n1206));
   DLY4X1 FE_PHC4795_n2015 (.Y(FE_PHN4795_n2015), 
	.A(n2015));
   DLY4X1 FE_PHC4794_n1636 (.Y(FE_PHN4794_n1636), 
	.A(n1636));
   DLY4X1 FE_PHC4793_n1357 (.Y(FE_PHN4793_n1357), 
	.A(n1357));
   DLY4X1 FE_PHC4792_n1643 (.Y(FE_PHN4792_n1643), 
	.A(n1643));
   DLY4X1 FE_PHC4791_n1550 (.Y(FE_PHN4791_n1550), 
	.A(n1550));
   DLY4X1 FE_PHC4790_n1237 (.Y(FE_PHN4790_n1237), 
	.A(n1237));
   DLY4X1 FE_PHC4789_n1053 (.Y(FE_PHN4789_n1053), 
	.A(n1053));
   DLY4X1 FE_PHC4788_n1912 (.Y(FE_PHN4788_n1912), 
	.A(n1912));
   DLY4X1 FE_PHC4787_n2314 (.Y(FE_PHN4787_n2314), 
	.A(n2314));
   DLY4X1 FE_PHC4786_n1922 (.Y(FE_PHN4786_n1922), 
	.A(n1922));
   DLY4X1 FE_PHC4785_n1150 (.Y(FE_PHN4785_n1150), 
	.A(n1150));
   DLY4X1 FE_PHC4784_n2022 (.Y(FE_PHN4784_n2022), 
	.A(n2022));
   DLY4X1 FE_PHC4783_n2383 (.Y(FE_PHN4783_n2383), 
	.A(n2383));
   DLY4X1 FE_PHC4782_n1164 (.Y(FE_PHN4782_n1164), 
	.A(n1164));
   DLY4X1 FE_PHC4781_n1605 (.Y(FE_PHN4781_n1605), 
	.A(n1605));
   DLY4X1 FE_PHC4780_n1294 (.Y(FE_PHN4780_n1294), 
	.A(n1294));
   DLY4X1 FE_PHC4779_n1987 (.Y(FE_PHN4779_n1987), 
	.A(n1987));
   DLY4X1 FE_PHC4778_n1043 (.Y(FE_PHN4778_n1043), 
	.A(n1043));
   DLY4X1 FE_PHC4777_n1103 (.Y(FE_PHN4777_n1103), 
	.A(n1103));
   DLY4X1 FE_PHC4776_n1651 (.Y(FE_PHN4776_n1651), 
	.A(n1651));
   DLY4X1 FE_PHC4775_n902 (.Y(FE_PHN4775_n902), 
	.A(n902));
   DLY4X1 FE_PHC4774_n1867 (.Y(FE_PHN4774_n1867), 
	.A(FE_PHN2689_n1867));
   DLY4X1 FE_PHC4773_n1980 (.Y(FE_PHN4773_n1980), 
	.A(n1980));
   DLY4X1 FE_PHC4772_n1638 (.Y(FE_PHN4772_n1638), 
	.A(n1638));
   DLY4X1 FE_PHC4771_n1529 (.Y(FE_PHN4771_n1529), 
	.A(n1529));
   DLY4X1 FE_PHC4770_n1078 (.Y(FE_PHN4770_n1078), 
	.A(n1078));
   DLY4X1 FE_PHC4769_n1129 (.Y(FE_PHN4769_n1129), 
	.A(n1129));
   DLY4X1 FE_PHC4768_n1615 (.Y(FE_PHN4768_n1615), 
	.A(n1615));
   DLY4X1 FE_PHC4767_n2369 (.Y(FE_PHN4767_n2369), 
	.A(n2369));
   DLY4X1 FE_PHC4766_n1213 (.Y(FE_PHN4766_n1213), 
	.A(n1213));
   DLY4X1 FE_PHC4765_n1157 (.Y(FE_PHN4765_n1157), 
	.A(n1157));
   DLY3X1 FE_PHC4764_n1177 (.Y(FE_PHN4764_n1177), 
	.A(n1177));
   DLY3X1 FE_PHC4763_n1302 (.Y(FE_PHN4763_n1302), 
	.A(n1302));
   DLY3X1 FE_PHC4762_n1059 (.Y(FE_PHN4762_n1059), 
	.A(n1059));
   DLY3X1 FE_PHC4761_n1276 (.Y(FE_PHN4761_n1276), 
	.A(n1276));
   DLY4X1 FE_PHC4760_n1564 (.Y(FE_PHN4760_n1564), 
	.A(n1564));
   DLY4X1 FE_PHC4759_n2024 (.Y(FE_PHN4759_n2024), 
	.A(n2024));
   DLY3X1 FE_PHC4758_n1202 (.Y(FE_PHN4758_n1202), 
	.A(n1202));
   DLY4X1 FE_PHC4757_n1216 (.Y(FE_PHN4757_n1216), 
	.A(n1216));
   DLY3X1 FE_PHC4756_n926 (.Y(FE_PHN4756_n926), 
	.A(n926));
   DLY4X1 FE_PHC4755_n1155 (.Y(FE_PHN4755_n1155), 
	.A(n1155));
   DLY4X1 FE_PHC4754_n1584 (.Y(FE_PHN4754_n1584), 
	.A(n1584));
   DLY4X1 FE_PHC4753_n1589 (.Y(FE_PHN4753_n1589), 
	.A(n1589));
   DLY4X1 FE_PHC4752_n1019 (.Y(FE_PHN4752_n1019), 
	.A(n1019));
   DLY4X1 FE_PHC4751_n920 (.Y(FE_PHN4751_n920), 
	.A(n920));
   DLY4X1 FE_PHC4750_n1200 (.Y(FE_PHN4750_n1200), 
	.A(n1200));
   DLY3X1 FE_PHC4749_n2114 (.Y(FE_PHN4749_n2114), 
	.A(FE_PHN2707_n2114));
   DLY4X1 FE_PHC4748_n1601 (.Y(FE_PHN4748_n1601), 
	.A(n1601));
   DLY4X1 FE_PHC4747_n2004 (.Y(FE_PHN4747_n2004), 
	.A(n2004));
   DLY4X1 FE_PHC4746_n1255 (.Y(FE_PHN4746_n1255), 
	.A(n1255));
   DLY4X1 FE_PHC4745_n1979 (.Y(FE_PHN4745_n1979), 
	.A(n1979));
   DLY4X1 FE_PHC4744_n1117 (.Y(FE_PHN4744_n1117), 
	.A(n1117));
   DLY4X1 FE_PHC4743_n1349 (.Y(FE_PHN4743_n1349), 
	.A(n1349));
   DLY4X1 FE_PHC4742_n1058 (.Y(FE_PHN4742_n1058), 
	.A(n1058));
   DLY4X1 FE_PHC4741_n1940 (.Y(FE_PHN4741_n1940), 
	.A(n1940));
   DLY4X1 FE_PHC4740_n1093 (.Y(FE_PHN4740_n1093), 
	.A(n1093));
   DLY4X1 FE_PHC4739_n1354 (.Y(FE_PHN4739_n1354), 
	.A(n1354));
   DLY4X1 FE_PHC4738_n1159 (.Y(FE_PHN4738_n1159), 
	.A(n1159));
   DLY4X1 FE_PHC4737_n1642 (.Y(FE_PHN4737_n1642), 
	.A(n1642));
   DLY4X1 FE_PHC4736_n1602 (.Y(FE_PHN4736_n1602), 
	.A(n1602));
   DLY4X1 FE_PHC4735_n1629 (.Y(FE_PHN4735_n1629), 
	.A(n1629));
   DLY4X1 FE_PHC4734_n2084 (.Y(FE_PHN4734_n2084), 
	.A(n2084));
   DLY4X1 FE_PHC4733_n1215 (.Y(FE_PHN4733_n1215), 
	.A(n1215));
   DLY4X1 FE_PHC4732_n973 (.Y(FE_PHN4732_n973), 
	.A(n973));
   DLY4X1 FE_PHC4731_n2188 (.Y(FE_PHN4731_n2188), 
	.A(n2188));
   DLY4X1 FE_PHC4730_n2180 (.Y(FE_PHN4730_n2180), 
	.A(n2180));
   DLY4X1 FE_PHC4729_n1935 (.Y(FE_PHN4729_n1935), 
	.A(n1935));
   DLY4X1 FE_PHC4728_n2033 (.Y(FE_PHN4728_n2033), 
	.A(n2033));
   DLY4X1 FE_PHC4727_n1338 (.Y(FE_PHN4727_n1338), 
	.A(n1338));
   DLY4X1 FE_PHC4726_n1195 (.Y(FE_PHN4726_n1195), 
	.A(n1195));
   DLY4X1 FE_PHC4725_n1138 (.Y(FE_PHN4725_n1138), 
	.A(n1138));
   DLY4X1 FE_PHC4724_n1365 (.Y(FE_PHN4724_n1365), 
	.A(n1365));
   DLY4X1 FE_PHC4723_n1167 (.Y(FE_PHN4723_n1167), 
	.A(n1167));
   DLY4X1 FE_PHC4722_n1990 (.Y(FE_PHN4722_n1990), 
	.A(n1990));
   DLY4X1 FE_PHC4721_n1887 (.Y(FE_PHN4721_n1887), 
	.A(n1887));
   DLY4X1 FE_PHC4720_n2256 (.Y(FE_PHN4720_n2256), 
	.A(n2256));
   DLY4X1 FE_PHC4719_n1075 (.Y(FE_PHN4719_n1075), 
	.A(n1075));
   DLY3X1 FE_PHC4718_n2209 (.Y(FE_PHN4718_n2209), 
	.A(n2209));
   DLY4X1 FE_PHC4717_n1110 (.Y(FE_PHN4717_n1110), 
	.A(n1110));
   DLY4X1 FE_PHC4716_n1622 (.Y(FE_PHN4716_n1622), 
	.A(n1622));
   DLY3X1 FE_PHC4715_n2320 (.Y(FE_PHN4715_n2320), 
	.A(n2320));
   DLY4X1 FE_PHC4714_n1284 (.Y(FE_PHN4714_n1284), 
	.A(n1284));
   DLY3X1 FE_PHC4713_n1283 (.Y(FE_PHN4713_n1283), 
	.A(n1283));
   DLY4X1 FE_PHC4712_n2031 (.Y(FE_PHN4712_n2031), 
	.A(n2031));
   DLY3X1 FE_PHC4711_n1640 (.Y(FE_PHN4711_n1640), 
	.A(n1640));
   DLY4X1 FE_PHC4710_n1131 (.Y(FE_PHN4710_n1131), 
	.A(n1131));
   DLY4X1 FE_PHC4709_n915 (.Y(FE_PHN4709_n915), 
	.A(n915));
   DLY4X1 FE_PHC4708_n1119 (.Y(FE_PHN4708_n1119), 
	.A(n1119));
   DLY3X1 FE_PHC4707_n1205 (.Y(FE_PHN4707_n1205), 
	.A(n1205));
   DLY4X1 FE_PHC4706_n1977 (.Y(FE_PHN4706_n1977), 
	.A(n1977));
   DLY3X1 FE_PHC4705_n2117 (.Y(FE_PHN4705_n2117), 
	.A(n2117));
   DLY4X1 FE_PHC4704_n1527 (.Y(FE_PHN4704_n1527), 
	.A(n1527));
   DLY4X1 FE_PHC4703_n2375 (.Y(FE_PHN4703_n2375), 
	.A(n2375));
   DLY4X1 FE_PHC4702_n1350 (.Y(FE_PHN4702_n1350), 
	.A(n1350));
   DLY3X1 FE_PHC4701_n2424 (.Y(FE_PHN4701_n2424), 
	.A(n2424));
   DLY4X1 FE_PHC4700_n1090 (.Y(FE_PHN4700_n1090), 
	.A(n1090));
   DLY4X1 FE_PHC4699_n1147 (.Y(FE_PHN4699_n1147), 
	.A(n1147));
   DLY3X1 FE_PHC4698_n1689 (.Y(FE_PHN4698_n1689), 
	.A(n1689));
   DLY4X1 FE_PHC4697_n1585 (.Y(FE_PHN4697_n1585), 
	.A(n1585));
   DLY3X1 FE_PHC4696_n953 (.Y(FE_PHN4696_n953), 
	.A(n953));
   DLY4X1 FE_PHC4695_n1949 (.Y(FE_PHN4695_n1949), 
	.A(n1949));
   DLY3X1 FE_PHC4694_n1125 (.Y(FE_PHN4694_n1125), 
	.A(n1125));
   DLY4X1 FE_PHC4693_n1944 (.Y(FE_PHN4693_n1944), 
	.A(n1944));
   DLY3X1 FE_PHC4692_n2201 (.Y(FE_PHN4692_n2201), 
	.A(n2201));
   DLY3X1 FE_PHC4691_n1929 (.Y(FE_PHN4691_n1929), 
	.A(n1929));
   DLY4X1 FE_PHC4690_n1641 (.Y(FE_PHN4690_n1641), 
	.A(n1641));
   DLY4X1 FE_PHC4689_n2030 (.Y(FE_PHN4689_n2030), 
	.A(n2030));
   DLY3X1 FE_PHC4688_n1551 (.Y(FE_PHN4688_n1551), 
	.A(n1551));
   DLY3X1 FE_PHC4687_n1339 (.Y(FE_PHN4687_n1339), 
	.A(n1339));
   DLY4X1 FE_PHC4686_n1183 (.Y(FE_PHN4686_n1183), 
	.A(n1183));
   DLY4X1 FE_PHC4685_n1528 (.Y(FE_PHN4685_n1528), 
	.A(n1528));
   DLY4X1 FE_PHC4684_n1746 (.Y(FE_PHN4684_n1746), 
	.A(n1746));
   DLY4X1 FE_PHC4683_n2011 (.Y(FE_PHN4683_n2011), 
	.A(n2011));
   DLY4X1 FE_PHC4682_n1392 (.Y(FE_PHN4682_n1392), 
	.A(n1392));
   DLY4X1 FE_PHC4681_n1533 (.Y(FE_PHN4681_n1533), 
	.A(n1533));
   DLY4X1 FE_PHC4680_n1130 (.Y(FE_PHN4680_n1130), 
	.A(n1130));
   DLY4X1 FE_PHC4679_n1553 (.Y(FE_PHN4679_n1553), 
	.A(n1553));
   DLY4X1 FE_PHC4678_n1303 (.Y(FE_PHN4678_n1303), 
	.A(n1303));
   DLY4X1 FE_PHC4677_n1098 (.Y(FE_PHN4677_n1098), 
	.A(n1098));
   DLY4X1 FE_PHC4676_n2060 (.Y(FE_PHN4676_n2060), 
	.A(n2060));
   DLY4X1 FE_PHC4675_n1992 (.Y(FE_PHN4675_n1992), 
	.A(n1992));
   DLY4X1 FE_PHC4674_n1315 (.Y(FE_PHN4674_n1315), 
	.A(n1315));
   DLY4X1 FE_PHC4673_n2330 (.Y(FE_PHN4673_n2330), 
	.A(n2330));
   DLY4X1 FE_PHC4672_n1235 (.Y(FE_PHN4672_n1235), 
	.A(n1235));
   DLY4X1 FE_PHC4671_n925 (.Y(FE_PHN4671_n925), 
	.A(n925));
   DLY4X1 FE_PHC4670_n1317 (.Y(FE_PHN4670_n1317), 
	.A(n1317));
   DLY4X1 FE_PHC4669_n1419 (.Y(FE_PHN4669_n1419), 
	.A(n1419));
   DLY4X1 FE_PHC4668_n1174 (.Y(FE_PHN4668_n1174), 
	.A(n1174));
   DLY4X1 FE_PHC4667_n1212 (.Y(FE_PHN4667_n1212), 
	.A(n1212));
   DLY4X1 FE_PHC4665_n2223 (.Y(FE_PHN4665_n2223), 
	.A(n2223));
   DLY4X1 FE_PHC4664_n2324 (.Y(FE_PHN4664_n2324), 
	.A(n2324));
   DLY4X1 FE_PHC4663_n1637 (.Y(FE_PHN4663_n1637), 
	.A(n1637));
   DLY4X1 FE_PHC4662_n936 (.Y(FE_PHN4662_n936), 
	.A(n936));
   DLY4X1 FE_PHC4661_n1324 (.Y(FE_PHN4661_n1324), 
	.A(n1324));
   DLY4X1 FE_PHC4660_n1322 (.Y(FE_PHN4660_n1322), 
	.A(n1322));
   DLY4X1 FE_PHC4659_n2016 (.Y(FE_PHN4659_n2016), 
	.A(n2016));
   DLY4X1 FE_PHC4658_n2305 (.Y(FE_PHN4658_n2305), 
	.A(n2305));
   DLY4X1 FE_PHC4657_n2116 (.Y(FE_PHN4657_n2116), 
	.A(n2116));
   DLY4X1 FE_PHC4656_n1226 (.Y(FE_PHN4656_n1226), 
	.A(n1226));
   DLY3X1 FE_PHC4655_n2081 (.Y(FE_PHN4655_n2081), 
	.A(n2081));
   DLY3X1 FE_PHC4654_n1610 (.Y(FE_PHN4654_n1610), 
	.A(n1610));
   DLY4X1 FE_PHC4653_n1069 (.Y(FE_PHN4653_n1069), 
	.A(n1069));
   DLY3X1 FE_PHC4652_n1959 (.Y(FE_PHN4652_n1959), 
	.A(n1959));
   DLY4X1 FE_PHC4651_n1566 (.Y(FE_PHN4651_n1566), 
	.A(n1566));
   DLY4X1 FE_PHC4650_n2316 (.Y(FE_PHN4650_n2316), 
	.A(n2316));
   DLY4X1 FE_PHC4649_n1108 (.Y(FE_PHN4649_n1108), 
	.A(n1108));
   DLY4X1 FE_PHC4648_n1025 (.Y(FE_PHN4648_n1025), 
	.A(n1025));
   DLY4X1 FE_PHC4647_n1036 (.Y(FE_PHN4647_n1036), 
	.A(n1036));
   DLY4X1 FE_PHC4646_n1188 (.Y(FE_PHN4646_n1188), 
	.A(n1188));
   DLY4X1 FE_PHC4644_n1532 (.Y(FE_PHN4644_n1532), 
	.A(n1532));
   DLY4X1 FE_PHC4643_n1352 (.Y(FE_PHN4643_n1352), 
	.A(n1352));
   DLY4X1 FE_PHC4642_n1569 (.Y(FE_PHN4642_n1569), 
	.A(n1569));
   DLY4X1 FE_PHC4641_n1363 (.Y(FE_PHN4641_n1363), 
	.A(n1363));
   DLY4X1 FE_PHC4640_n1120 (.Y(FE_PHN4640_n1120), 
	.A(n1120));
   DLY4X1 FE_PHC4639_n1145 (.Y(FE_PHN4639_n1145), 
	.A(n1145));
   DLY3X1 FE_PHC4638_n1123 (.Y(FE_PHN4638_n1123), 
	.A(n1123));
   DLY4X1 FE_PHC4637_n1219 (.Y(FE_PHN4637_n1219), 
	.A(n1219));
   DLY3X1 FE_PHC4636_n1321 (.Y(FE_PHN4636_n1321), 
	.A(n1321));
   DLY3X1 FE_PHC4635_n1613 (.Y(FE_PHN4635_n1613), 
	.A(n1613));
   DLY4X1 FE_PHC4634_n2119 (.Y(FE_PHN4634_n2119), 
	.A(n2119));
   DLY4X1 FE_PHC4633_n1538 (.Y(FE_PHN4633_n1538), 
	.A(n1538));
   DLY3X1 FE_PHC4632_n1915 (.Y(FE_PHN4632_n1915), 
	.A(n1915));
   DLY3X1 FE_PHC4631_n2275 (.Y(FE_PHN4631_n2275), 
	.A(n2275));
   DLY3X1 FE_PHC4630_n1575 (.Y(FE_PHN4630_n1575), 
	.A(n1575));
   DLY3X1 FE_PHC4629_n2368 (.Y(FE_PHN4629_n2368), 
	.A(n2368));
   DLY3X1 FE_PHC4628_n932 (.Y(FE_PHN4628_n932), 
	.A(n932));
   DLY4X1 FE_PHC4627_n1072 (.Y(FE_PHN4627_n1072), 
	.A(n1072));
   DLY4X1 FE_PHC4626_n1272 (.Y(FE_PHN4626_n1272), 
	.A(n1272));
   DLY4X1 FE_PHC4625_n1570 (.Y(FE_PHN4625_n1570), 
	.A(n1570));
   DLY4X1 FE_PHC4624_n1556 (.Y(FE_PHN4624_n1556), 
	.A(n1556));
   DLY4X1 FE_PHC4623_n1836 (.Y(FE_PHN4623_n1836), 
	.A(n1836));
   DLY3X1 FE_PHC4622_n1806 (.Y(FE_PHN4622_n1806), 
	.A(n1806));
   DLY4X1 FE_PHC4621_n1924 (.Y(FE_PHN4621_n1924), 
	.A(n1924));
   DLY4X1 FE_PHC4620_n1313 (.Y(FE_PHN4620_n1313), 
	.A(n1313));
   DLY4X1 FE_PHC4619_n1026 (.Y(FE_PHN4619_n1026), 
	.A(n1026));
   DLY4X1 FE_PHC4618_n1007 (.Y(FE_PHN4618_n1007), 
	.A(n1007));
   DLY4X1 FE_PHC4617_n2014 (.Y(FE_PHN4617_n2014), 
	.A(n2014));
   DLY3X1 FE_PHC4616_n2155 (.Y(FE_PHN4616_n2155), 
	.A(n2155));
   DLY3X1 FE_PHC4615_n1281 (.Y(FE_PHN4615_n1281), 
	.A(n1281));
   DLY3X1 FE_PHC4614_n907 (.Y(FE_PHN4614_n907), 
	.A(n907));
   DLY3X1 FE_PHC4613_n1583 (.Y(FE_PHN4613_n1583), 
	.A(n1583));
   DLY4X1 FE_PHC4612_n887 (.Y(FE_PHN4612_n887), 
	.A(n887));
   DLY4X1 FE_PHC4611_n1525 (.Y(FE_PHN4611_n1525), 
	.A(n1525));
   DLY4X1 FE_PHC4610_n1133 (.Y(FE_PHN4610_n1133), 
	.A(n1133));
   DLY4X1 FE_PHC4609_n2019 (.Y(FE_PHN4609_n2019), 
	.A(n2019));
   DLY3X1 FE_PHC4608_n2283 (.Y(FE_PHN4608_n2283), 
	.A(n2283));
   DLY3X1 FE_PHC4607_n909 (.Y(FE_PHN4607_n909), 
	.A(n909));
   DLY4X1 FE_PHC4606_n1381 (.Y(FE_PHN4606_n1381), 
	.A(n1381));
   DLY4X1 FE_PHC4605_n1176 (.Y(FE_PHN4605_n1176), 
	.A(n1176));
   DLY4X1 FE_PHC4604_n1136 (.Y(FE_PHN4604_n1136), 
	.A(n1136));
   DLY4X1 FE_PHC4603_n2139 (.Y(FE_PHN4603_n2139), 
	.A(n2139));
   DLY4X1 FE_PHC4602_n1548 (.Y(FE_PHN4602_n1548), 
	.A(n1548));
   DLY4X1 FE_PHC4601_n1972 (.Y(FE_PHN4601_n1972), 
	.A(n1972));
   DLY4X1 FE_PHC4600_n1182 (.Y(FE_PHN4600_n1182), 
	.A(n1182));
   DLY4X1 FE_PHC4599_n1380 (.Y(FE_PHN4599_n1380), 
	.A(n1380));
   DLY4X1 FE_PHC4598_n1582 (.Y(FE_PHN4598_n1582), 
	.A(n1582));
   DLY4X1 FE_PHC4597_n960 (.Y(FE_PHN4597_n960), 
	.A(n960));
   DLY4X1 FE_PHC4596_n977 (.Y(FE_PHN4596_n977), 
	.A(n977));
   DLY4X1 FE_PHC4595_n1388 (.Y(FE_PHN4595_n1388), 
	.A(n1388));
   DLY4X1 FE_PHC4594_n1934 (.Y(FE_PHN4594_n1934), 
	.A(n1934));
   DLY4X1 FE_PHC4593_n1387 (.Y(FE_PHN4593_n1387), 
	.A(n1387));
   DLY4X1 FE_PHC4592_n1543 (.Y(FE_PHN4592_n1543), 
	.A(n1543));
   DLY4X1 FE_PHC4591_n2310 (.Y(FE_PHN4591_n2310), 
	.A(n2310));
   DLY4X1 FE_PHC4590_n1332 (.Y(FE_PHN4590_n1332), 
	.A(n1332));
   DLY4X1 FE_PHC4589_n948 (.Y(FE_PHN4589_n948), 
	.A(n948));
   DLY4X1 FE_PHC4588_n2049 (.Y(FE_PHN4588_n2049), 
	.A(n2049));
   DLY4X1 FE_PHC4587_n1744 (.Y(FE_PHN4587_n1744), 
	.A(FE_PHN2747_n1744));
   DLY4X1 FE_PHC4586_n1918 (.Y(FE_PHN4586_n1918), 
	.A(n1918));
   DLY4X1 FE_PHC4585_n1970 (.Y(FE_PHN4585_n1970), 
	.A(n1970));
   DLY4X1 FE_PHC4584_n1986 (.Y(FE_PHN4584_n1986), 
	.A(n1986));
   DLY4X1 FE_PHC4583_n1211 (.Y(FE_PHN4583_n1211), 
	.A(n1211));
   DLY4X1 FE_PHC4582_n1982 (.Y(FE_PHN4582_n1982), 
	.A(n1982));
   DLY4X1 FE_PHC4581_n1623 (.Y(FE_PHN4581_n1623), 
	.A(n1623));
   DLY4X1 FE_PHC4580_n1857 (.Y(FE_PHN4580_n1857), 
	.A(n1857));
   DLY4X1 FE_PHC4579_n1018 (.Y(FE_PHN4579_n1018), 
	.A(n1018));
   DLY4X1 FE_PHC4578_n1068 (.Y(FE_PHN4578_n1068), 
	.A(n1068));
   DLY4X1 FE_PHC4577_n1812 (.Y(FE_PHN4577_n1812), 
	.A(n1812));
   DLY4X1 FE_PHC4576_n1092 (.Y(FE_PHN4576_n1092), 
	.A(n1092));
   DLY4X1 FE_PHC4575_n2309 (.Y(FE_PHN4575_n2309), 
	.A(n2309));
   DLY4X1 FE_PHC4574_n1639 (.Y(FE_PHN4574_n1639), 
	.A(n1639));
   DLY4X1 FE_PHC4573_n1015 (.Y(FE_PHN4573_n1015), 
	.A(n1015));
   DLY4X1 FE_PHC4572_n2005 (.Y(FE_PHN4572_n2005), 
	.A(n2005));
   DLY4X1 FE_PHC4571_n1914 (.Y(FE_PHN4571_n1914), 
	.A(n1914));
   DLY3X1 FE_PHC4570_n2007 (.Y(FE_PHN4570_n2007), 
	.A(n2007));
   DLY4X1 FE_PHC4569_n1132 (.Y(FE_PHN4569_n1132), 
	.A(n1132));
   DLY4X1 FE_PHC4568_n1331 (.Y(FE_PHN4568_n1331), 
	.A(n1331));
   DLY4X1 FE_PHC4567_n2185 (.Y(FE_PHN4567_n2185), 
	.A(n2185));
   DLY4X1 FE_PHC4566_n1952 (.Y(FE_PHN4566_n1952), 
	.A(n1952));
   DLY3X1 FE_PHC4565_n1820 (.Y(FE_PHN4565_n1820), 
	.A(n1820));
   DLY4X1 FE_PHC4564_n2384 (.Y(FE_PHN4564_n2384), 
	.A(n2384));
   DLY4X1 FE_PHC4563_n1966 (.Y(FE_PHN4563_n1966), 
	.A(n1966));
   DLY4X1 FE_PHC4562_n2010 (.Y(FE_PHN4562_n2010), 
	.A(n2010));
   DLY4X1 FE_PHC4561_n1044 (.Y(FE_PHN4561_n1044), 
	.A(n1044));
   DLY4X1 FE_PHC4560_n1383 (.Y(FE_PHN4560_n1383), 
	.A(n1383));
   DLY4X1 FE_PHC4559_n1190 (.Y(FE_PHN4559_n1190), 
	.A(n1190));
   DLY3X1 FE_PHC4558_n1947 (.Y(FE_PHN4558_n1947), 
	.A(n1947));
   DLY4X1 FE_PHC4557_n1181 (.Y(FE_PHN4557_n1181), 
	.A(n1181));
   DLY4X1 FE_PHC4556_n1005 (.Y(FE_PHN4556_n1005), 
	.A(n1005));
   DLY4X1 FE_PHC4555_n1245 (.Y(FE_PHN4555_n1245), 
	.A(n1245));
   DLY4X1 FE_PHC4554_n999 (.Y(FE_PHN4554_n999), 
	.A(n999));
   DLY4X1 FE_PHC4553_n1113 (.Y(FE_PHN4553_n1113), 
	.A(n1113));
   DLY4X1 FE_PHC4552_n1360 (.Y(FE_PHN4552_n1360), 
	.A(n1360));
   DLY3X1 FE_PHC4551_n1579 (.Y(FE_PHN4551_n1579), 
	.A(n1579));
   DLY4X1 FE_PHC4550_n1559 (.Y(FE_PHN4550_n1559), 
	.A(n1559));
   DLY4X1 FE_PHC4549_n1361 (.Y(FE_PHN4549_n1361), 
	.A(n1361));
   DLY4X1 FE_PHC4548_n1534 (.Y(FE_PHN4548_n1534), 
	.A(n1534));
   DLY3X1 FE_PHC4547_n2182 (.Y(FE_PHN4547_n2182), 
	.A(n2182));
   DLY4X1 FE_PHC4546_n1080 (.Y(FE_PHN4546_n1080), 
	.A(n1080));
   DLY4X1 FE_PHC4545_n1146 (.Y(FE_PHN4545_n1146), 
	.A(n1146));
   DLY3X1 FE_PHC4544_n1004 (.Y(FE_PHN4544_n1004), 
	.A(n1004));
   DLY3X1 FE_PHC4543_n1006 (.Y(FE_PHN4543_n1006), 
	.A(n1006));
   DLY4X1 FE_PHC4542_n2046 (.Y(FE_PHN4542_n2046), 
	.A(FE_PHN2693_n2046));
   DLY4X1 FE_PHC4541_n1187 (.Y(FE_PHN4541_n1187), 
	.A(n1187));
   DLY4X1 FE_PHC4540_n1050 (.Y(FE_PHN4540_n1050), 
	.A(n1050));
   DLY4X1 FE_PHC4539_n1057 (.Y(FE_PHN4539_n1057), 
	.A(n1057));
   DLY4X1 FE_PHC4538_n1034 (.Y(FE_PHN4538_n1034), 
	.A(n1034));
   DLY4X1 FE_PHC4537_n2094 (.Y(FE_PHN4537_n2094), 
	.A(n2094));
   DLY4X1 FE_PHC4536_n2307 (.Y(FE_PHN4536_n2307), 
	.A(n2307));
   DLY4X1 FE_PHC4535_n1358 (.Y(FE_PHN4535_n1358), 
	.A(n1358));
   DLY4X1 FE_PHC4534_n1229 (.Y(FE_PHN4534_n1229), 
	.A(n1229));
   DLY4X1 FE_PHC4533_n1151 (.Y(FE_PHN4533_n1151), 
	.A(n1151));
   DLY3X1 FE_PHC4532_n1552 (.Y(FE_PHN4532_n1552), 
	.A(n1552));
   DLY3X1 FE_PHC4531_n1650 (.Y(FE_PHN4531_n1650), 
	.A(n1650));
   DLY4X1 FE_PHC4530_n2388 (.Y(FE_PHN4530_n2388), 
	.A(n2388));
   DLY3X1 FE_PHC4529_n1462 (.Y(FE_PHN4529_n1462), 
	.A(n1462));
   DLY4X1 FE_PHC4528_n1135 (.Y(FE_PHN4528_n1135), 
	.A(n1135));
   DLY4X1 FE_PHC4527_n1562 (.Y(FE_PHN4527_n1562), 
	.A(n1562));
   DLY4X1 FE_PHC4526_n2191 (.Y(FE_PHN4526_n2191), 
	.A(n2191));
   DLY3X1 FE_PHC4525_n943 (.Y(FE_PHN4525_n943), 
	.A(n943));
   DLY4X1 FE_PHC4524_n1826 (.Y(FE_PHN4524_n1826), 
	.A(n1826));
   DLY4X1 FE_PHC4523_n1035 (.Y(FE_PHN4523_n1035), 
	.A(n1035));
   DLY4X1 FE_PHC4522_n1049 (.Y(FE_PHN4522_n1049), 
	.A(n1049));
   DLY3X1 FE_PHC4521_n1386 (.Y(FE_PHN4521_n1386), 
	.A(n1386));
   DLY4X1 FE_PHC4520_n1101 (.Y(FE_PHN4520_n1101), 
	.A(n1101));
   DLY4X1 FE_PHC4519_n1345 (.Y(FE_PHN4519_n1345), 
	.A(n1345));
   DLY3X1 FE_PHC4518_n1985 (.Y(FE_PHN4518_n1985), 
	.A(n1985));
   DLY4X1 FE_PHC4517_n1879 (.Y(FE_PHN4517_n1879), 
	.A(n1879));
   DLY3X1 FE_PHC4516_n1624 (.Y(FE_PHN4516_n1624), 
	.A(n1624));
   DLY4X1 FE_PHC4515_n1379 (.Y(FE_PHN4515_n1379), 
	.A(n1379));
   DLY4X1 FE_PHC4514_n1493 (.Y(FE_PHN4514_n1493), 
	.A(FE_PHN2671_n1493));
   DLY4X1 FE_PHC4513_n1728 (.Y(FE_PHN4513_n1728), 
	.A(n1728));
   DLY4X1 FE_PHC4512_n1170 (.Y(FE_PHN4512_n1170), 
	.A(n1170));
   DLY4X1 FE_PHC4511_n1468 (.Y(FE_PHN4511_n1468), 
	.A(n1468));
   DLY4X1 FE_PHC4510_n1341 (.Y(FE_PHN4510_n1341), 
	.A(n1341));
   DLY4X1 FE_PHC4509_n1201 (.Y(FE_PHN4509_n1201), 
	.A(n1201));
   DLY4X1 FE_PHC4508_n1163 (.Y(FE_PHN4508_n1163), 
	.A(n1163));
   DLY4X1 FE_PHC4507_n1169 (.Y(FE_PHN4507_n1169), 
	.A(n1169));
   DLY4X1 FE_PHC4506_n1153 (.Y(FE_PHN4506_n1153), 
	.A(n1153));
   DLY4X1 FE_PHC4505_n1936 (.Y(FE_PHN4505_n1936), 
	.A(n1936));
   DLY4X1 FE_PHC4504_n1652 (.Y(FE_PHN4504_n1652), 
	.A(n1652));
   DLY4X1 FE_PHC4503_n1278 (.Y(FE_PHN4503_n1278), 
	.A(n1278));
   DLY4X1 FE_PHC4502_n1755 (.Y(FE_PHN4502_n1755), 
	.A(n1755));
   DLY4X1 FE_PHC4501_n1084 (.Y(FE_PHN4501_n1084), 
	.A(n1084));
   DLY4X1 FE_PHC4500_n1197 (.Y(FE_PHN4500_n1197), 
	.A(n1197));
   DLY4X1 FE_PHC4499_n1008 (.Y(FE_PHN4499_n1008), 
	.A(n1008));
   DLY4X1 FE_PHC4498_n1731 (.Y(FE_PHN4498_n1731), 
	.A(n1731));
   DLY4X1 FE_PHC4497_n1950 (.Y(FE_PHN4497_n1950), 
	.A(n1950));
   DLY4X1 FE_PHC4496_n912 (.Y(FE_PHN4496_n912), 
	.A(n912));
   DLY4X1 FE_PHC4495_n1046 (.Y(FE_PHN4495_n1046), 
	.A(n1046));
   DLY4X1 FE_PHC4494_n914 (.Y(FE_PHN4494_n914), 
	.A(n914));
   DLY4X1 FE_PHC4493_n1376 (.Y(FE_PHN4493_n1376), 
	.A(n1376));
   DLY4X1 FE_PHC4492_n1572 (.Y(FE_PHN4492_n1572), 
	.A(n1572));
   DLY4X1 FE_PHC4491_n1974 (.Y(FE_PHN4491_n1974), 
	.A(n1974));
   DLY4X1 FE_PHC4490_n1925 (.Y(FE_PHN4490_n1925), 
	.A(n1925));
   DLY4X1 FE_PHC4489_n2311 (.Y(FE_PHN4489_n2311), 
	.A(n2311));
   DLY4X1 FE_PHC4488_n1910 (.Y(FE_PHN4488_n1910), 
	.A(n1910));
   DLY4X1 FE_PHC4487_n2159 (.Y(FE_PHN4487_n2159), 
	.A(n2159));
   DLY4X1 FE_PHC4486_n1536 (.Y(FE_PHN4486_n1536), 
	.A(n1536));
   DLY4X1 FE_PHC4485_n1234 (.Y(FE_PHN4485_n1234), 
	.A(n1234));
   DLY4X1 FE_PHC4484_n1061 (.Y(FE_PHN4484_n1061), 
	.A(n1061));
   DLY4X1 FE_PHC4483_n928 (.Y(FE_PHN4483_n928), 
	.A(n928));
   DLY4X1 FE_PHC4482_n1325 (.Y(FE_PHN4482_n1325), 
	.A(n1325));
   DLY4X1 FE_PHC4481_n927 (.Y(FE_PHN4481_n927), 
	.A(n927));
   DLY4X1 FE_PHC4480_n1988 (.Y(FE_PHN4480_n1988), 
	.A(n1988));
   DLY4X1 FE_PHC4479_n2238 (.Y(FE_PHN4479_n2238), 
	.A(n2238));
   DLY4X1 FE_PHC4478_n1688 (.Y(FE_PHN4478_n1688), 
	.A(n1688));
   DLY4X1 FE_PHC4477_n2301 (.Y(FE_PHN4477_n2301), 
	.A(n2301));
   DLY4X1 FE_PHC4476_n1779 (.Y(FE_PHN4476_n1779), 
	.A(n1779));
   DLY4X1 FE_PHC4475_n1865 (.Y(FE_PHN4475_n1865), 
	.A(n1865));
   DLY4X1 FE_PHC4474_n1645 (.Y(FE_PHN4474_n1645), 
	.A(n1645));
   DLY4X1 FE_PHC4473_n1312 (.Y(FE_PHN4473_n1312), 
	.A(n1312));
   DLY3X1 FE_PHC4472_n1856 (.Y(FE_PHN4472_n1856), 
	.A(n1856));
   DLY4X1 FE_PHC4471_n1089 (.Y(FE_PHN4471_n1089), 
	.A(n1089));
   DLY3X1 FE_PHC4470_n1031 (.Y(FE_PHN4470_n1031), 
	.A(n1031));
   DLY4X1 FE_PHC4469_n1592 (.Y(FE_PHN4469_n1592), 
	.A(n1592));
   DLY4X1 FE_PHC4468_n1942 (.Y(FE_PHN4468_n1942), 
	.A(n1942));
   DLY3X1 FE_PHC4467_n896 (.Y(FE_PHN4467_n896), 
	.A(n896));
   DLY4X1 FE_PHC4466_n942 (.Y(FE_PHN4466_n942), 
	.A(n942));
   DLY4X1 FE_PHC4465_n1014 (.Y(FE_PHN4465_n1014), 
	.A(n1014));
   DLY4X1 FE_PHC4464_n1634 (.Y(FE_PHN4464_n1634), 
	.A(n1634));
   DLY4X1 FE_PHC4463_n1628 (.Y(FE_PHN4463_n1628), 
	.A(n1628));
   DLY4X1 FE_PHC4462_n2382 (.Y(FE_PHN4462_n2382), 
	.A(n2382));
   DLY3X1 FE_PHC4461_n1514 (.Y(FE_PHN4461_n1514), 
	.A(n1514));
   DLY4X1 FE_PHC4460_n1083 (.Y(FE_PHN4460_n1083), 
	.A(n1083));
   DLY4X1 FE_PHC4459_n1993 (.Y(FE_PHN4459_n1993), 
	.A(n1993));
   DLY3X1 FE_PHC4458_n2138 (.Y(FE_PHN4458_n2138), 
	.A(n2138));
   DLY4X1 FE_PHC4457_n2322 (.Y(FE_PHN4457_n2322), 
	.A(n2322));
   DLY4X1 FE_PHC4456_n1384 (.Y(FE_PHN4456_n1384), 
	.A(n1384));
   DLY3X1 FE_PHC4455_n1588 (.Y(FE_PHN4455_n1588), 
	.A(n1588));
   DLY4X1 FE_PHC4454_n1270 (.Y(FE_PHN4454_n1270), 
	.A(n1270));
   DLY4X1 FE_PHC4453_n1122 (.Y(FE_PHN4453_n1122), 
	.A(n1122));
   DLY3X1 FE_PHC4452_n2228 (.Y(FE_PHN4452_n2228), 
	.A(FE_PHN2670_n2228));
   DLY3X1 FE_PHC4451_n1683 (.Y(FE_PHN4451_n1683), 
	.A(n1683));
   DLY3X1 FE_PHC4450_n2167 (.Y(FE_PHN4450_n2167), 
	.A(n2167));
   DLY3X1 FE_PHC4449_n2149 (.Y(FE_PHN4449_n2149), 
	.A(n2149));
   DLY4X1 FE_PHC4448_n2325 (.Y(FE_PHN4448_n2325), 
	.A(n2325));
   DLY3X1 FE_PHC4447_n1047 (.Y(FE_PHN4447_n1047), 
	.A(n1047));
   DLY3X1 FE_PHC4446_n1595 (.Y(FE_PHN4446_n1595), 
	.A(FE_PHN1812_n1595));
   DLY3X1 FE_PHC4445_n1635 (.Y(FE_PHN4445_n1635), 
	.A(n1635));
   DLY4X1 FE_PHC4444_n1927 (.Y(FE_PHN4444_n1927), 
	.A(n1927));
   DLY4X1 FE_PHC4443_n1568 (.Y(FE_PHN4443_n1568), 
	.A(n1568));
   DLY4X1 FE_PHC4442_n2148 (.Y(FE_PHN4442_n2148), 
	.A(n2148));
   DLY4X1 FE_PHC4441_n1269 (.Y(FE_PHN4441_n1269), 
	.A(n1269));
   DLY3X1 FE_PHC4440_n1832 (.Y(FE_PHN4440_n1832), 
	.A(n1832));
   DLY4X1 FE_PHC4439_n1076 (.Y(FE_PHN4439_n1076), 
	.A(n1076));
   DLY4X1 FE_PHC4438_n1260 (.Y(FE_PHN4438_n1260), 
	.A(n1260));
   DLY4X1 FE_PHC4437_n1969 (.Y(FE_PHN4437_n1969), 
	.A(n1969));
   DLY4X1 FE_PHC4436_n1625 (.Y(FE_PHN4436_n1625), 
	.A(n1625));
   DLY3X1 FE_PHC4435_n2232 (.Y(FE_PHN4435_n2232), 
	.A(n2232));
   DLY4X1 FE_PHC4434_n1401 (.Y(FE_PHN4434_n1401), 
	.A(n1401));
   DLY3X1 FE_PHC4433_n1373 (.Y(FE_PHN4433_n1373), 
	.A(n1373));
   DLY4X1 FE_PHC4432_n1168 (.Y(FE_PHN4432_n1168), 
	.A(n1168));
   DLY4X1 FE_PHC4431_n1295 (.Y(FE_PHN4431_n1295), 
	.A(n1295));
   DLY4X1 FE_PHC4430_n945 (.Y(FE_PHN4430_n945), 
	.A(n945));
   DLY4X1 FE_PHC4429_n1343 (.Y(FE_PHN4429_n1343), 
	.A(n1343));
   DLY4X1 FE_PHC4428_n1432 (.Y(FE_PHN4428_n1432), 
	.A(n1432));
   DLY3X1 FE_PHC4427_n1813 (.Y(FE_PHN4427_n1813), 
	.A(n1813));
   DLY4X1 FE_PHC4426_n1540 (.Y(FE_PHN4426_n1540), 
	.A(n1540));
   DLY4X1 FE_PHC4425_n1242 (.Y(FE_PHN4425_n1242), 
	.A(n1242));
   DLY4X1 FE_PHC4424_n1166 (.Y(FE_PHN4424_n1166), 
	.A(n1166));
   DLY4X1 FE_PHC4423_n1378 (.Y(FE_PHN4423_n1378), 
	.A(n1378));
   DLY4X1 FE_PHC4422_n1971 (.Y(FE_PHN4422_n1971), 
	.A(n1971));
   DLY4X1 FE_PHC4421_n2009 (.Y(FE_PHN4421_n2009), 
	.A(n2009));
   DLY4X1 FE_PHC4420_n1853 (.Y(FE_PHN4420_n1853), 
	.A(n1853));
   DLY4X1 FE_PHC4419_n1734 (.Y(FE_PHN4419_n1734), 
	.A(n1734));
   DLY4X1 FE_PHC4418_n1056 (.Y(FE_PHN4418_n1056), 
	.A(n1056));
   DLY4X1 FE_PHC4417_n2378 (.Y(FE_PHN4417_n2378), 
	.A(n2378));
   DLY4X1 FE_PHC4416_n1286 (.Y(FE_PHN4416_n1286), 
	.A(n1286));
   DLY4X1 FE_PHC4415_n1374 (.Y(FE_PHN4415_n1374), 
	.A(n1374));
   DLY4X1 FE_PHC4414_n1094 (.Y(FE_PHN4414_n1094), 
	.A(n1094));
   DLY4X1 FE_PHC4413_n1064 (.Y(FE_PHN4413_n1064), 
	.A(n1064));
   DLY4X1 FE_PHC4412_n2306 (.Y(FE_PHN4412_n2306), 
	.A(n2306));
   DLY4X1 FE_PHC4411_n1960 (.Y(FE_PHN4411_n1960), 
	.A(n1960));
   DLY4X1 FE_PHC4410_n1955 (.Y(FE_PHN4410_n1955), 
	.A(n1955));
   DLY4X1 FE_PHC4409_n956 (.Y(FE_PHN4409_n956), 
	.A(n956));
   DLY4X1 FE_PHC4408_n2234 (.Y(FE_PHN4408_n2234), 
	.A(n2234));
   DLY4X1 FE_PHC4407_n1573 (.Y(FE_PHN4407_n1573), 
	.A(n1573));
   DLY4X1 FE_PHC4406_n1838 (.Y(FE_PHN4406_n1838), 
	.A(n1838));
   DLY4X1 FE_PHC4405_n1298 (.Y(FE_PHN4405_n1298), 
	.A(n1298));
   DLY4X1 FE_PHC4404_n921 (.Y(FE_PHN4404_n921), 
	.A(n921));
   DLY4X1 FE_PHC4403_n1051 (.Y(FE_PHN4403_n1051), 
	.A(n1051));
   DLY4X1 FE_PHC4402_n1603 (.Y(FE_PHN4402_n1603), 
	.A(n1603));
   DLY4X1 FE_PHC4401_n1218 (.Y(FE_PHN4401_n1218), 
	.A(n1218));
   DLY4X1 FE_PHC4400_n1140 (.Y(FE_PHN4400_n1140), 
	.A(n1140));
   DLY4X1 FE_PHC4399_n1554 (.Y(FE_PHN4399_n1554), 
	.A(n1554));
   DLY4X1 FE_PHC4398_n1368 (.Y(FE_PHN4398_n1368), 
	.A(n1368));
   DLY4X1 FE_PHC4397_n2321 (.Y(FE_PHN4397_n2321), 
	.A(n2321));
   DLY4X1 FE_PHC4396_n2387 (.Y(FE_PHN4396_n2387), 
	.A(n2387));
   DLY4X1 FE_PHC4395_n983 (.Y(FE_PHN4395_n983), 
	.A(n983));
   DLY4X1 FE_PHC4394_n1535 (.Y(FE_PHN4394_n1535), 
	.A(n1535));
   DLY4X1 FE_PHC4393_n2267 (.Y(FE_PHN4393_n2267), 
	.A(n2267));
   DLY4X1 FE_PHC4392_n1917 (.Y(FE_PHN4392_n1917), 
	.A(n1917));
   DLY4X1 FE_PHC4391_n1265 (.Y(FE_PHN4391_n1265), 
	.A(n1265));
   DLY4X1 FE_PHC4390_n1292 (.Y(FE_PHN4390_n1292), 
	.A(n1292));
   DLY4X1 FE_PHC4389_n1478 (.Y(FE_PHN4389_n1478), 
	.A(n1478));
   DLY4X1 FE_PHC4388_n1956 (.Y(FE_PHN4388_n1956), 
	.A(n1956));
   DLY4X1 FE_PHC4387_n1530 (.Y(FE_PHN4387_n1530), 
	.A(n1530));
   DLY4X1 FE_PHC4386_n1749 (.Y(FE_PHN4386_n1749), 
	.A(n1749));
   DLY4X1 FE_PHC4385_n1892 (.Y(FE_PHN4385_n1892), 
	.A(n1892));
   DLY4X1 FE_PHC4384_n2194 (.Y(FE_PHN4384_n2194), 
	.A(n2194));
   DLY4X1 FE_PHC4383_n1288 (.Y(FE_PHN4383_n1288), 
	.A(n1288));
   DLY4X1 FE_PHC4382_n963 (.Y(FE_PHN4382_n963), 
	.A(n963));
   DLY4X1 FE_PHC4381_n1184 (.Y(FE_PHN4381_n1184), 
	.A(n1184));
   DLY3X1 FE_PHC4380_n1464 (.Y(FE_PHN4380_n1464), 
	.A(n1464));
   DLY3X1 FE_PHC4379_n1758 (.Y(FE_PHN4379_n1758), 
	.A(FE_PHN2638_n1758));
   DLY4X1 FE_PHC4378_n1776 (.Y(FE_PHN4378_n1776), 
	.A(n1776));
   DLY3X1 FE_PHC4377_n1644 (.Y(FE_PHN4377_n1644), 
	.A(n1644));
   DLY3X1 FE_PHC4376_n1767 (.Y(FE_PHN4376_n1767), 
	.A(n1767));
   DLY4X1 FE_PHC4375_n2018 (.Y(FE_PHN4375_n2018), 
	.A(n2018));
   DLY4X1 FE_PHC4374_n1160 (.Y(FE_PHN4374_n1160), 
	.A(n1160));
   DLY4X1 FE_PHC4373_n1289 (.Y(FE_PHN4373_n1289), 
	.A(n1289));
   DLY3X1 FE_PHC4372_n1217 (.Y(FE_PHN4372_n1217), 
	.A(n1217));
   DLY3X1 FE_PHC4371_n1287 (.Y(FE_PHN4371_n1287), 
	.A(n1287));
   DLY4X1 FE_PHC4370_n998 (.Y(FE_PHN4370_n998), 
	.A(n998));
   DLY3X1 FE_PHC4369_n1240 (.Y(FE_PHN4369_n1240), 
	.A(n1240));
   DLY4X1 FE_PHC4368_n1077 (.Y(FE_PHN4368_n1077), 
	.A(n1077));
   DLY4X1 FE_PHC4367_n1097 (.Y(FE_PHN4367_n1097), 
	.A(n1097));
   DLY4X1 FE_PHC4366_n1028 (.Y(FE_PHN4366_n1028), 
	.A(n1028));
   DLY4X1 FE_PHC4365_n1953 (.Y(FE_PHN4365_n1953), 
	.A(n1953));
   DLY4X1 FE_PHC4364_n1391 (.Y(FE_PHN4364_n1391), 
	.A(n1391));
   DLY4X1 FE_PHC4363_n1351 (.Y(FE_PHN4363_n1351), 
	.A(n1351));
   DLY4X1 FE_PHC4362_n1227 (.Y(FE_PHN4362_n1227), 
	.A(n1227));
   DLY4X1 FE_PHC4361_n1377 (.Y(FE_PHN4361_n1377), 
	.A(n1377));
   DLY4X1 FE_PHC4360_n1810 (.Y(FE_PHN4360_n1810), 
	.A(n1810));
   DLY4X1 FE_PHC4359_n2174 (.Y(FE_PHN4359_n2174), 
	.A(n2174));
   DLY3X1 FE_PHC4358_n2157 (.Y(FE_PHN4358_n2157), 
	.A(n2157));
   DLY4X1 FE_PHC4357_n1016 (.Y(FE_PHN4357_n1016), 
	.A(n1016));
   DLY4X1 FE_PHC4356_n1306 (.Y(FE_PHN4356_n1306), 
	.A(n1306));
   DLY4X1 FE_PHC4355_n1675 (.Y(FE_PHN4355_n1675), 
	.A(n1675));
   DLY4X1 FE_PHC4354_n1908 (.Y(FE_PHN4354_n1908), 
	.A(n1908));
   DLY4X1 FE_PHC4353_n1697 (.Y(FE_PHN4353_n1697), 
	.A(n1697));
   DLY3X1 FE_PHC4352_n1296 (.Y(FE_PHN4352_n1296), 
	.A(n1296));
   DLY4X1 FE_PHC4351_n1366 (.Y(FE_PHN4351_n1366), 
	.A(n1366));
   DLY4X1 FE_PHC4350_n1105 (.Y(FE_PHN4350_n1105), 
	.A(n1105));
   DLY4X1 FE_PHC4349_n1560 (.Y(FE_PHN4349_n1560), 
	.A(n1560));
   DLY4X1 FE_PHC4348_n2020 (.Y(FE_PHN4348_n2020), 
	.A(n2020));
   DLY4X1 FE_PHC4347_n1861 (.Y(FE_PHN4347_n1861), 
	.A(n1861));
   DLY4X1 FE_PHC4346_n2008 (.Y(FE_PHN4346_n2008), 
	.A(n2008));
   DLY4X1 FE_PHC4345_n1964 (.Y(FE_PHN4345_n1964), 
	.A(n1964));
   DLY4X1 FE_PHC4344_n1479 (.Y(FE_PHN4344_n1479), 
	.A(n1479));
   DLY4X1 FE_PHC4343_n1342 (.Y(FE_PHN4343_n1342), 
	.A(n1342));
   DLY4X1 FE_PHC4342_n1695 (.Y(FE_PHN4342_n1695), 
	.A(n1695));
   DLY3X1 FE_PHC4341_n1275 (.Y(FE_PHN4341_n1275), 
	.A(n1275));
   DLY4X1 FE_PHC4340_n1414 (.Y(FE_PHN4340_n1414), 
	.A(n1414));
   DLY4X1 FE_PHC4339_n1946 (.Y(FE_PHN4339_n1946), 
	.A(n1946));
   DLY4X1 FE_PHC4338_n1938 (.Y(FE_PHN4338_n1938), 
	.A(n1938));
   DLY4X1 FE_PHC4337_n1238 (.Y(FE_PHN4337_n1238), 
	.A(n1238));
   DLY4X1 FE_PHC4336_n975 (.Y(FE_PHN4336_n975), 
	.A(n975));
   DLY4X1 FE_PHC4335_n1843 (.Y(FE_PHN4335_n1843), 
	.A(FE_PHN2617_n1843));
   DLY4X1 FE_PHC4334_n1461 (.Y(FE_PHN4334_n1461), 
	.A(n1461));
   DLY4X1 FE_PHC4333_n2317 (.Y(FE_PHN4333_n2317), 
	.A(n2317));
   DLY4X1 FE_PHC4332_n1670 (.Y(FE_PHN4332_n1670), 
	.A(n1670));
   DLY4X1 FE_PHC4331_n2253 (.Y(FE_PHN4331_n2253), 
	.A(n2253));
   DLY4X1 FE_PHC4330_n1791 (.Y(FE_PHN4330_n1791), 
	.A(n1791));
   DLY4X1 FE_PHC4329_n2023 (.Y(FE_PHN4329_n2023), 
	.A(n2023));
   DLY4X1 FE_PHC4328_n1060 (.Y(FE_PHN4328_n1060), 
	.A(n1060));
   DLY4X1 FE_PHC4327_n1505 (.Y(FE_PHN4327_n1505), 
	.A(n1505));
   DLY4X1 FE_PHC4326_n1633 (.Y(FE_PHN4326_n1633), 
	.A(n1633));
   DLY4X1 FE_PHC4325_n929 (.Y(FE_PHN4325_n929), 
	.A(n929));
   DLY4X1 FE_PHC4324_n1372 (.Y(FE_PHN4324_n1372), 
	.A(n1372));
   DLY4X1 FE_PHC4323_n1859 (.Y(FE_PHN4323_n1859), 
	.A(n1859));
   DLY4X1 FE_PHC4322_n2025 (.Y(FE_PHN4322_n2025), 
	.A(n2025));
   DLY4X1 FE_PHC4321_n1301 (.Y(FE_PHN4321_n1301), 
	.A(n1301));
   DLY4X1 FE_PHC4320_n1079 (.Y(FE_PHN4320_n1079), 
	.A(n1079));
   DLY4X1 FE_PHC4319_n961 (.Y(FE_PHN4319_n961), 
	.A(n961));
   DLY4X1 FE_PHC4318_n1396 (.Y(FE_PHN4318_n1396), 
	.A(n1396));
   DLY4X1 FE_PHC4317_n1340 (.Y(FE_PHN4317_n1340), 
	.A(n1340));
   DLY4X1 FE_PHC4316_n978 (.Y(FE_PHN4316_n978), 
	.A(n978));
   DLY4X1 FE_PHC4315_n1305 (.Y(FE_PHN4315_n1305), 
	.A(n1305));
   DLY4X1 FE_PHC4314_n1663 (.Y(FE_PHN4314_n1663), 
	.A(n1663));
   DLY4X1 FE_PHC4313_n1648 (.Y(FE_PHN4313_n1648), 
	.A(n1648));
   DLY4X1 FE_PHC4312_n1968 (.Y(FE_PHN4312_n1968), 
	.A(n1968));
   DLY4X1 FE_PHC4311_n1096 (.Y(FE_PHN4311_n1096), 
	.A(n1096));
   DLY4X1 FE_PHC4310_n1225 (.Y(FE_PHN4310_n1225), 
	.A(n1225));
   DLY4X1 FE_PHC4309_n1346 (.Y(FE_PHN4309_n1346), 
	.A(n1346));
   DLY4X1 FE_PHC4308_n1362 (.Y(FE_PHN4308_n1362), 
	.A(n1362));
   DLY4X1 FE_PHC4307_n1104 (.Y(FE_PHN4307_n1104), 
	.A(n1104));
   DLY4X1 FE_PHC4306_n1389 (.Y(FE_PHN4306_n1389), 
	.A(n1389));
   DLY4X1 FE_PHC4305_n2013 (.Y(FE_PHN4305_n2013), 
	.A(n2013));
   DLY4X1 FE_PHC4304_n2328 (.Y(FE_PHN4304_n2328), 
	.A(n2328));
   DLY4X1 FE_PHC4303_n900 (.Y(FE_PHN4303_n900), 
	.A(n900));
   DLY4X1 FE_PHC4302_n947 (.Y(FE_PHN4302_n947), 
	.A(n947));
   DLY4X1 FE_PHC4301_n1222 (.Y(FE_PHN4301_n1222), 
	.A(n1222));
   DLY4X1 FE_PHC4300_n1477 (.Y(FE_PHN4300_n1477), 
	.A(n1477));
   DLY4X1 FE_PHC4299_n2029 (.Y(FE_PHN4299_n2029), 
	.A(n2029));
   DLY4X1 FE_PHC4298_n2172 (.Y(FE_PHN4298_n2172), 
	.A(n2172));
   DLY4X1 FE_PHC4297_n2258 (.Y(FE_PHN4297_n2258), 
	.A(n2258));
   DLY4X1 FE_PHC4296_n1074 (.Y(FE_PHN4296_n1074), 
	.A(n1074));
   DLY4X1 FE_PHC4295_n1082 (.Y(FE_PHN4295_n1082), 
	.A(n1082));
   DLY4X1 FE_PHC4294_n976 (.Y(FE_PHN4294_n976), 
	.A(n976));
   DLY4X1 FE_PHC4293_n1790 (.Y(FE_PHN4293_n1790), 
	.A(n1790));
   DLY4X1 FE_PHC4292_n2027 (.Y(FE_PHN4292_n2027), 
	.A(n2027));
   DLY4X1 FE_PHC4291_n1591 (.Y(FE_PHN4291_n1591), 
	.A(n1591));
   DLY4X1 FE_PHC4290_n1845 (.Y(FE_PHN4290_n1845), 
	.A(n1845));
   DLY4X1 FE_PHC4289_n1926 (.Y(FE_PHN4289_n1926), 
	.A(n1926));
   DLY4X1 FE_PHC4288_n1700 (.Y(FE_PHN4288_n1700), 
	.A(n1700));
   DLY4X1 FE_PHC4287_n1042 (.Y(FE_PHN4287_n1042), 
	.A(n1042));
   DLY4X1 FE_PHC4286_n1280 (.Y(FE_PHN4286_n1280), 
	.A(n1280));
   DLY4X1 FE_PHC4285_n2380 (.Y(FE_PHN4285_n2380), 
	.A(n2380));
   DLY4X1 FE_PHC4284_n2065 (.Y(FE_PHN4284_n2065), 
	.A(n2065));
   DLY4X1 FE_PHC4283_n1654 (.Y(FE_PHN4283_n1654), 
	.A(n1654));
   DLY4X1 FE_PHC4282_n1816 (.Y(FE_PHN4282_n1816), 
	.A(n1816));
   DLY3X1 FE_PHC4281_n1291 (.Y(FE_PHN4281_n1291), 
	.A(n1291));
   DLY4X1 FE_PHC4280_n2239 (.Y(FE_PHN4280_n2239), 
	.A(n2239));
   DLY4X1 FE_PHC4279_n2156 (.Y(FE_PHN4279_n2156), 
	.A(n2156));
   DLY3X1 FE_PHC4278_n1963 (.Y(FE_PHN4278_n1963), 
	.A(n1963));
   DLY4X1 FE_PHC4277_n916 (.Y(FE_PHN4277_n916), 
	.A(n916));
   DLY4X1 FE_PHC4276_n1277 (.Y(FE_PHN4276_n1277), 
	.A(n1277));
   DLY3X1 FE_PHC4275_n1279 (.Y(FE_PHN4275_n1279), 
	.A(n1279));
   DLY4X1 FE_PHC4274_n2271 (.Y(FE_PHN4274_n2271), 
	.A(n2271));
   DLY4X1 FE_PHC4273_n2111 (.Y(FE_PHN4273_n2111), 
	.A(n2111));
   DLY4X1 FE_PHC4272_n2026 (.Y(FE_PHN4272_n2026), 
	.A(n2026));
   DLY4X1 FE_PHC4271_n1931 (.Y(FE_PHN4271_n1931), 
	.A(n1931));
   DLY4X1 FE_PHC4270_n1930 (.Y(FE_PHN4270_n1930), 
	.A(n1930));
   DLY3X1 FE_PHC4269_n2323 (.Y(FE_PHN4269_n2323), 
	.A(n2323));
   DLY4X1 FE_PHC4268_n1567 (.Y(FE_PHN4268_n1567), 
	.A(n1567));
   DLY4X1 FE_PHC4267_n2115 (.Y(FE_PHN4267_n2115), 
	.A(n2115));
   DLY4X1 FE_PHC4266_n2226 (.Y(FE_PHN4266_n2226), 
	.A(n2226));
   DLY4X1 FE_PHC4265_n1496 (.Y(FE_PHN4265_n1496), 
	.A(n1496));
   DLY4X1 FE_PHC4264_n1983 (.Y(FE_PHN4264_n1983), 
	.A(n1983));
   DLY3X1 FE_PHC4263_n2329 (.Y(FE_PHN4263_n2329), 
	.A(n2329));
   DLY4X1 FE_PHC4262_n1107 (.Y(FE_PHN4262_n1107), 
	.A(n1107));
   DLY4X1 FE_PHC4261_n1991 (.Y(FE_PHN4261_n1991), 
	.A(n1991));
   DLY4X1 FE_PHC4260_n2179 (.Y(FE_PHN4260_n2179), 
	.A(n2179));
   DLY4X1 FE_PHC4259_n2140 (.Y(FE_PHN4259_n2140), 
	.A(n2140));
   DLY4X1 FE_PHC4258_n2032 (.Y(FE_PHN4258_n2032), 
	.A(n2032));
   DLY4X1 FE_PHC4257_n2207 (.Y(FE_PHN4257_n2207), 
	.A(n2207));
   DLY4X1 FE_PHC4256_n934 (.Y(FE_PHN4256_n934), 
	.A(n934));
   DLY4X1 FE_PHC4255_n1911 (.Y(FE_PHN4255_n1911), 
	.A(n1911));
   DLY4X1 FE_PHC4254_n2184 (.Y(FE_PHN4254_n2184), 
	.A(n2184));
   DLY4X1 FE_PHC4253_n1102 (.Y(FE_PHN4253_n1102), 
	.A(n1102));
   DLY4X1 FE_PHC4252_n1081 (.Y(FE_PHN4252_n1081), 
	.A(n1081));
   DLY4X1 FE_PHC4251_n1484 (.Y(FE_PHN4251_n1484), 
	.A(n1484));
   DLY4X1 FE_PHC4250_n1881 (.Y(FE_PHN4250_n1881), 
	.A(n1881));
   DLY4X1 FE_PHC4249_n1748 (.Y(FE_PHN4249_n1748), 
	.A(n1748));
   DLY4X1 FE_PHC4248_n2012 (.Y(FE_PHN4248_n2012), 
	.A(n2012));
   DLY4X1 FE_PHC4247_n1370 (.Y(FE_PHN4247_n1370), 
	.A(n1370));
   DLY4X1 FE_PHC4246_n1017 (.Y(FE_PHN4246_n1017), 
	.A(n1017));
   DLY4X1 FE_PHC4245_n1954 (.Y(FE_PHN4245_n1954), 
	.A(n1954));
   DLY4X1 FE_PHC4244_n1445 (.Y(FE_PHN4244_n1445), 
	.A(n1445));
   DLY3X1 FE_PHC4243_n1909 (.Y(FE_PHN4243_n1909), 
	.A(n1909));
   DLY4X1 FE_PHC4242_n2280 (.Y(FE_PHN4242_n2280), 
	.A(n2280));
   DLY4X1 FE_PHC4241_n1347 (.Y(FE_PHN4241_n1347), 
	.A(n1347));
   DLY4X1 FE_PHC4240_n1236 (.Y(FE_PHN4240_n1236), 
	.A(n1236));
   DLY4X1 FE_PHC4239_n1112 (.Y(FE_PHN4239_n1112), 
	.A(n1112));
   DLY4X1 FE_PHC4238_n1784 (.Y(FE_PHN4238_n1784), 
	.A(n1784));
   DLY4X1 FE_PHC4237_n1839 (.Y(FE_PHN4237_n1839), 
	.A(n1839));
   DLY4X1 FE_PHC4236_n2045 (.Y(FE_PHN4236_n2045), 
	.A(n2045));
   DLY4X1 FE_PHC4235_n1825 (.Y(FE_PHN4235_n1825), 
	.A(n1825));
   DLY4X1 FE_PHC4234_n1054 (.Y(FE_PHN4234_n1054), 
	.A(n1054));
   DLY4X1 FE_PHC4233_n952 (.Y(FE_PHN4233_n952), 
	.A(n952));
   DLY4X1 FE_PHC4232_n1480 (.Y(FE_PHN4232_n1480), 
	.A(n1480));
   DLY4X1 FE_PHC4231_n1574 (.Y(FE_PHN4231_n1574), 
	.A(n1574));
   DLY4X1 FE_PHC4230_n1783 (.Y(FE_PHN4230_n1783), 
	.A(n1783));
   DLY4X1 FE_PHC4229_n959 (.Y(FE_PHN4229_n959), 
	.A(n959));
   DLY4X1 FE_PHC4228_n1765 (.Y(FE_PHN4228_n1765), 
	.A(n1765));
   DLY4X1 FE_PHC4227_n1961 (.Y(FE_PHN4227_n1961), 
	.A(n1961));
   DLY4X1 FE_PHC4226_n1040 (.Y(FE_PHN4226_n1040), 
	.A(n1040));
   DLY4X1 FE_PHC4225_n1609 (.Y(FE_PHN4225_n1609), 
	.A(n1609));
   DLY4X1 FE_PHC4224_n1707 (.Y(FE_PHN4224_n1707), 
	.A(n1707));
   DLY4X1 FE_PHC4223_n1735 (.Y(FE_PHN4223_n1735), 
	.A(n1735));
   DLY4X1 FE_PHC4222_n913 (.Y(FE_PHN4222_n913), 
	.A(n913));
   DLY4X1 FE_PHC4221_n1780 (.Y(FE_PHN4221_n1780), 
	.A(n1780));
   DLY4X1 FE_PHC4220_n2061 (.Y(FE_PHN4220_n2061), 
	.A(n2061));
   DLY4X1 FE_PHC4219_n1590 (.Y(FE_PHN4219_n1590), 
	.A(n1590));
   DLY4X1 FE_PHC4218_n1830 (.Y(FE_PHN4218_n1830), 
	.A(n1830));
   DLY4X1 FE_PHC4217_n1257 (.Y(FE_PHN4217_n1257), 
	.A(n1257));
   DLY4X1 FE_PHC4216_n1111 (.Y(FE_PHN4216_n1111), 
	.A(n1111));
   DLY4X1 FE_PHC4215_n2189 (.Y(FE_PHN4215_n2189), 
	.A(FE_PHN2645_n2189));
   DLY4X1 FE_PHC4214_n1516 (.Y(FE_PHN4214_n1516), 
	.A(n1516));
   DLY4X1 FE_PHC4213_n919 (.Y(FE_PHN4213_n919), 
	.A(n919));
   DLY4X1 FE_PHC4212_n911 (.Y(FE_PHN4212_n911), 
	.A(n911));
   DLY4X1 FE_PHC4211_n1510 (.Y(FE_PHN4211_n1510), 
	.A(n1510));
   DLY4X1 FE_PHC4210_n1996 (.Y(FE_PHN4210_n1996), 
	.A(n1996));
   DLY4X1 FE_PHC4209_n2123 (.Y(FE_PHN4209_n2123), 
	.A(n2123));
   DLY4X1 FE_PHC4208_n1385 (.Y(FE_PHN4208_n1385), 
	.A(n1385));
   DLY4X1 FE_PHC4207_n1995 (.Y(FE_PHN4207_n1995), 
	.A(n1995));
   DLY4X1 FE_PHC4206_n2047 (.Y(FE_PHN4206_n2047), 
	.A(n2047));
   DLY4X1 FE_PHC4205_n1841 (.Y(FE_PHN4205_n1841), 
	.A(n1841));
   DLY4X1 FE_PHC4204_n1024 (.Y(FE_PHN4204_n1024), 
	.A(n1024));
   DLY4X1 FE_PHC4203_n2151 (.Y(FE_PHN4203_n2151), 
	.A(n2151));
   DLY4X1 FE_PHC4202_n2071 (.Y(FE_PHN4202_n2071), 
	.A(n2071));
   DLY4X1 FE_PHC4201_n1751 (.Y(FE_PHN4201_n1751), 
	.A(n1751));
   DLY4X1 FE_PHC4200_n1620 (.Y(FE_PHN4200_n1620), 
	.A(n1620));
   DLY4X1 FE_PHC4199_n1837 (.Y(FE_PHN4199_n1837), 
	.A(n1837));
   DLY4X1 FE_PHC4198_n1766 (.Y(FE_PHN4198_n1766), 
	.A(n1766));
   DLY4X1 FE_PHC4197_n1668 (.Y(FE_PHN4197_n1668), 
	.A(n1668));
   DLY4X1 FE_PHC4196_n2144 (.Y(FE_PHN4196_n2144), 
	.A(n2144));
   DLY4X1 FE_PHC4195_n2318 (.Y(FE_PHN4195_n2318), 
	.A(n2318));
   DLY4X1 FE_PHC4194_n1520 (.Y(FE_PHN4194_n1520), 
	.A(n1520));
   DLY4X1 FE_PHC4193_n2052 (.Y(FE_PHN4193_n2052), 
	.A(n2052));
   DLY4X1 FE_PHC4192_n970 (.Y(FE_PHN4192_n970), 
	.A(n970));
   DLY4X1 FE_PHC4191_n1032 (.Y(FE_PHN4191_n1032), 
	.A(n1032));
   DLY4X1 FE_PHC4190_n1885 (.Y(FE_PHN4190_n1885), 
	.A(n1885));
   DLY4X1 FE_PHC4189_n2367 (.Y(FE_PHN4189_n2367), 
	.A(n2367));
   DLY4X1 FE_PHC4188_n1828 (.Y(FE_PHN4188_n1828), 
	.A(n1828));
   DLY4X1 FE_PHC4187_n1063 (.Y(FE_PHN4187_n1063), 
	.A(n1063));
   DLY4X1 FE_PHC4186_n1418 (.Y(FE_PHN4186_n1418), 
	.A(n1418));
   DLY4X1 FE_PHC4185_n1311 (.Y(FE_PHN4185_n1311), 
	.A(n1311));
   DLY4X1 FE_PHC4184_n2287 (.Y(FE_PHN4184_n2287), 
	.A(FE_PHN2604_n2287));
   DLY4X1 FE_PHC4183_n1541 (.Y(FE_PHN4183_n1541), 
	.A(n1541));
   DLY4X1 FE_PHC4182_n1407 (.Y(FE_PHN4182_n1407), 
	.A(n1407));
   DLY4X1 FE_PHC4181_n1375 (.Y(FE_PHN4181_n1375), 
	.A(n1375));
   DLY4X1 FE_PHC4180_n2038 (.Y(FE_PHN4180_n2038), 
	.A(n2038));
   DLY4X1 FE_PHC4179_n2278 (.Y(FE_PHN4179_n2278), 
	.A(n2278));
   DLY4X1 FE_PHC4178_n1504 (.Y(FE_PHN4178_n1504), 
	.A(n1504));
   DLY4X1 FE_PHC4177_n1831 (.Y(FE_PHN4177_n1831), 
	.A(n1831));
   DLY4X1 FE_PHC4176_n1250 (.Y(FE_PHN4176_n1250), 
	.A(n1250));
   DLY4X1 FE_PHC4175_n1430 (.Y(FE_PHN4175_n1430), 
	.A(n1430));
   DLY4X1 FE_PHC4174_n1455 (.Y(FE_PHN4174_n1455), 
	.A(n1455));
   DLY4X1 FE_PHC4173_n1676 (.Y(FE_PHN4173_n1676), 
	.A(n1676));
   DLY4X1 FE_PHC4172_n2040 (.Y(FE_PHN4172_n2040), 
	.A(n2040));
   DLY4X1 FE_PHC4171_n1507 (.Y(FE_PHN4171_n1507), 
	.A(n1507));
   DLY4X1 FE_PHC4170_n1161 (.Y(FE_PHN4170_n1161), 
	.A(n1161));
   DLY4X1 FE_PHC4169_n2093 (.Y(FE_PHN4169_n2093), 
	.A(n2093));
   DLY4X1 FE_PHC4168_n1958 (.Y(FE_PHN4168_n1958), 
	.A(n1958));
   DLY4X1 FE_PHC4167_n1808 (.Y(FE_PHN4167_n1808), 
	.A(n1808));
   DLY4X1 FE_PHC4166_n2163 (.Y(FE_PHN4166_n2163), 
	.A(n2163));
   DLY4X1 FE_PHC4165_n1309 (.Y(FE_PHN4165_n1309), 
	.A(n1309));
   DLY4X1 FE_PHC4164_n1124 (.Y(FE_PHN4164_n1124), 
	.A(n1124));
   DLY4X1 FE_PHC4163_n2043 (.Y(FE_PHN4163_n2043), 
	.A(n2043));
   DLY4X1 FE_PHC4162_n1742 (.Y(FE_PHN4162_n1742), 
	.A(n1742));
   DLY4X1 FE_PHC4161_n1409 (.Y(FE_PHN4161_n1409), 
	.A(n1409));
   DLY4X1 FE_PHC4160_n1420 (.Y(FE_PHN4160_n1420), 
	.A(n1420));
   DLY4X1 FE_PHC4159_n1427 (.Y(FE_PHN4159_n1427), 
	.A(n1427));
   DLY4X1 FE_PHC4158_n2222 (.Y(FE_PHN4158_n2222), 
	.A(n2222));
   DLY4X1 FE_PHC4157_n1500 (.Y(FE_PHN4157_n1500), 
	.A(n1500));
   DLY4X1 FE_PHC4156_n2241 (.Y(FE_PHN4156_n2241), 
	.A(n2241));
   DLY4X1 FE_PHC4155_n2064 (.Y(FE_PHN4155_n2064), 
	.A(n2064));
   DLY4X1 FE_PHC4154_n1937 (.Y(FE_PHN4154_n1937), 
	.A(n1937));
   DLY4X1 FE_PHC4153_n1565 (.Y(FE_PHN4153_n1565), 
	.A(n1565));
   DLY4X1 FE_PHC4152_n1545 (.Y(FE_PHN4152_n1545), 
	.A(n1545));
   DLY4X1 FE_PHC4151_n1335 (.Y(FE_PHN4151_n1335), 
	.A(n1335));
   DLY4X1 FE_PHC4150_n1330 (.Y(FE_PHN4150_n1330), 
	.A(n1330));
   DLY4X1 FE_PHC4149_n1011 (.Y(FE_PHN4149_n1011), 
	.A(n1011));
   DLY4X1 FE_PHC4148_n1677 (.Y(FE_PHN4148_n1677), 
	.A(n1677));
   DLY4X1 FE_PHC4147_n979 (.Y(FE_PHN4147_n979), 
	.A(n979));
   DLY4X1 FE_PHC4146_n933 (.Y(FE_PHN4146_n933), 
	.A(n933));
   DLY4X1 FE_PHC4145_n1299 (.Y(FE_PHN4145_n1299), 
	.A(n1299));
   DLY4X1 FE_PHC4144_n1900 (.Y(FE_PHN4144_n1900), 
	.A(n1900));
   DLY4X1 FE_PHC4143_n1799 (.Y(FE_PHN4143_n1799), 
	.A(n1799));
   DLY4X1 FE_PHC4142_n1449 (.Y(FE_PHN4142_n1449), 
	.A(n1449));
   DLY4X1 FE_PHC4141_n1410 (.Y(FE_PHN4141_n1410), 
	.A(n1410));
   DLY4X1 FE_PHC4140_n2147 (.Y(FE_PHN4140_n2147), 
	.A(n2147));
   DLY4X1 FE_PHC4139_n971 (.Y(FE_PHN4139_n971), 
	.A(n971));
   DLY4X1 FE_PHC4138_n1903 (.Y(FE_PHN4138_n1903), 
	.A(n1903));
   DLY4X1 FE_PHC4137_n1320 (.Y(FE_PHN4137_n1320), 
	.A(n1320));
   DLY4X1 FE_PHC4136_n1071 (.Y(FE_PHN4136_n1071), 
	.A(n1071));
   DLY4X1 FE_PHC4135_n2289 (.Y(FE_PHN4135_n2289), 
	.A(n2289));
   DLY4X1 FE_PHC4134_n984 (.Y(FE_PHN4134_n984), 
	.A(n984));
   DLY4X1 FE_PHC4133_n2216 (.Y(FE_PHN4133_n2216), 
	.A(n2216));
   DLY4X1 FE_PHC4132_n1665 (.Y(FE_PHN4132_n1665), 
	.A(n1665));
   DLY4X1 FE_PHC4131_n1907 (.Y(FE_PHN4131_n1907), 
	.A(n1907));
   DLY4X1 FE_PHC4130_n2131 (.Y(FE_PHN4130_n2131), 
	.A(n2131));
   DLY4X1 FE_PHC4129_n1088 (.Y(FE_PHN4129_n1088), 
	.A(n1088));
   DLY4X1 FE_PHC4128_n888 (.Y(FE_PHN4128_n888), 
	.A(n888));
   DLY4X1 FE_PHC4127_n940 (.Y(FE_PHN4127_n940), 
	.A(n940));
   DLY4X1 FE_PHC4126_n904 (.Y(FE_PHN4126_n904), 
	.A(n904));
   DLY4X1 FE_PHC4125_n937 (.Y(FE_PHN4125_n937), 
	.A(n937));
   DLY4X1 FE_PHC4124_n895 (.Y(FE_PHN4124_n895), 
	.A(n895));
   DLY4X1 FE_PHC4123_n1773 (.Y(FE_PHN4123_n1773), 
	.A(n1773));
   DLY4X1 FE_PHC4122_n1518 (.Y(FE_PHN4122_n1518), 
	.A(n1518));
   DLY4X1 FE_PHC4121_n1851 (.Y(FE_PHN4121_n1851), 
	.A(n1851));
   DLY4X1 FE_PHC4120_n2153 (.Y(FE_PHN4120_n2153), 
	.A(n2153));
   DLY4X1 FE_PHC4119_n1716 (.Y(FE_PHN4119_n1716), 
	.A(n1716));
   DLY4X1 FE_PHC4118_n2377 (.Y(FE_PHN4118_n2377), 
	.A(n2377));
   DLY4X1 FE_PHC4117_n2303 (.Y(FE_PHN4117_n2303), 
	.A(n2303));
   DLY4X1 FE_PHC4116_n1127 (.Y(FE_PHN4116_n1127), 
	.A(n1127));
   DLY4X1 FE_PHC4115_n1254 (.Y(FE_PHN4115_n1254), 
	.A(n1254));
   DLY4X1 FE_PHC4114_n1775 (.Y(FE_PHN4114_n1775), 
	.A(n1775));
   DLY4X1 FE_PHC4113_n1469 (.Y(FE_PHN4113_n1469), 
	.A(n1469));
   DLY4X1 FE_PHC4112_n1457 (.Y(FE_PHN4112_n1457), 
	.A(n1457));
   DLY4X1 FE_PHC4111_n1923 (.Y(FE_PHN4111_n1923), 
	.A(n1923));
   DLY4X1 FE_PHC4110_n1884 (.Y(FE_PHN4110_n1884), 
	.A(n1884));
   DLY4X1 FE_PHC4109_n1777 (.Y(FE_PHN4109_n1777), 
	.A(n1777));
   DLY4X1 FE_PHC4108_n1353 (.Y(FE_PHN4108_n1353), 
	.A(n1353));
   DLY4X1 FE_PHC4107_n1782 (.Y(FE_PHN4107_n1782), 
	.A(n1782));
   DLY4X1 FE_PHC4106_n2164 (.Y(FE_PHN4106_n2164), 
	.A(n2164));
   DLY4X1 FE_PHC4105_n1788 (.Y(FE_PHN4105_n1788), 
	.A(n1788));
   DLY4X1 FE_PHC4104_n1485 (.Y(FE_PHN4104_n1485), 
	.A(n1485));
   DLY4X1 FE_PHC4103_n1337 (.Y(FE_PHN4103_n1337), 
	.A(n1337));
   DLY4X1 FE_PHC4102_n1095 (.Y(FE_PHN4102_n1095), 
	.A(n1095));
   DLY4X1 FE_PHC4101_n2248 (.Y(FE_PHN4101_n2248), 
	.A(n2248));
   DLY3X1 FE_PHC4100_n1616 (.Y(FE_PHN4100_n1616), 
	.A(n1616));
   DLY4X1 FE_PHC4099_n2128 (.Y(FE_PHN4099_n2128), 
	.A(n2128));
   DLY4X1 FE_PHC4098_n1627 (.Y(FE_PHN4098_n1627), 
	.A(n1627));
   DLY4X1 FE_PHC4097_n2331 (.Y(FE_PHN4097_n2331), 
	.A(n2331));
   DLY4X1 FE_PHC4096_n1273 (.Y(FE_PHN4096_n1273), 
	.A(n1273));
   DLY4X1 FE_PHC4095_n2039 (.Y(FE_PHN4095_n2039), 
	.A(n2039));
   DLY4X1 FE_PHC4094_n1435 (.Y(FE_PHN4094_n1435), 
	.A(n1435));
   DLY4X1 FE_PHC4093_n1606 (.Y(FE_PHN4093_n1606), 
	.A(n1606));
   DLY4X1 FE_PHC4092_n1951 (.Y(FE_PHN4092_n1951), 
	.A(n1951));
   DLY4X1 FE_PHC4091_n2291 (.Y(FE_PHN4091_n2291), 
	.A(n2291));
   DLY4X1 FE_PHC4090_n1318 (.Y(FE_PHN4090_n1318), 
	.A(n1318));
   DLY4X1 FE_PHC4089_n1513 (.Y(FE_PHN4089_n1513), 
	.A(n1513));
   DLY4X1 FE_PHC4088_n2021 (.Y(FE_PHN4088_n2021), 
	.A(n2021));
   DLY4X1 FE_PHC4087_n1333 (.Y(FE_PHN4087_n1333), 
	.A(n1333));
   DLY4X1 FE_PHC4086_n1708 (.Y(FE_PHN4086_n1708), 
	.A(n1708));
   DLY3X1 FE_PHC4085_n1471 (.Y(FE_PHN4085_n1471), 
	.A(n1471));
   DLY4X1 FE_PHC4084_n1659 (.Y(FE_PHN4084_n1659), 
	.A(n1659));
   DLY4X1 FE_PHC4083_n1920 (.Y(FE_PHN4083_n1920), 
	.A(n1920));
   DLY4X1 FE_PHC4082_n1626 (.Y(FE_PHN4082_n1626), 
	.A(n1626));
   DLY4X1 FE_PHC4081_n2236 (.Y(FE_PHN4081_n2236), 
	.A(n2236));
   DLY4X1 FE_PHC4080_n1271 (.Y(FE_PHN4080_n1271), 
	.A(n1271));
   DLY4X1 FE_PHC4079_n1336 (.Y(FE_PHN4079_n1336), 
	.A(n1336));
   DLY4X1 FE_PHC4078_n2292 (.Y(FE_PHN4078_n2292), 
	.A(n2292));
   DLY4X1 FE_PHC4077_n2240 (.Y(FE_PHN4077_n2240), 
	.A(n2240));
   DLY4X1 FE_PHC4076_n1862 (.Y(FE_PHN4076_n1862), 
	.A(n1862));
   DLY4X1 FE_PHC4075_n2003 (.Y(FE_PHN4075_n2003), 
	.A(n2003));
   DLY4X1 FE_PHC4074_n968 (.Y(FE_PHN4074_n968), 
	.A(n968));
   DLY4X1 FE_PHC4073_n1274 (.Y(FE_PHN4073_n1274), 
	.A(n1274));
   DLY4X1 FE_PHC4072_n1196 (.Y(FE_PHN4072_n1196), 
	.A(n1196));
   DLY3X1 FE_PHC4071_n1770 (.Y(FE_PHN4071_n1770), 
	.A(n1770));
   DLY4X1 FE_PHC4070_n1792 (.Y(FE_PHN4070_n1792), 
	.A(n1792));
   DLY4X1 FE_PHC4069_n1899 (.Y(FE_PHN4069_n1899), 
	.A(n1899));
   DLY4X1 FE_PHC4068_n1334 (.Y(FE_PHN4068_n1334), 
	.A(n1334));
   DLY4X1 FE_PHC4067_n2176 (.Y(FE_PHN4067_n2176), 
	.A(n2176));
   DLY4X1 FE_PHC4066_n2002 (.Y(FE_PHN4066_n2002), 
	.A(n2002));
   DLY4X1 FE_PHC4065_n1997 (.Y(FE_PHN4065_n1997), 
	.A(n1997));
   DLY4X1 FE_PHC4064_n1736 (.Y(FE_PHN4064_n1736), 
	.A(n1736));
   DLY4X1 FE_PHC4063_n2090 (.Y(FE_PHN4063_n2090), 
	.A(n2090));
   DLY4X1 FE_PHC4062_n1975 (.Y(FE_PHN4062_n1975), 
	.A(n1975));
   DLY4X1 FE_PHC4061_n1542 (.Y(FE_PHN4061_n1542), 
	.A(n1542));
   DLY4X1 FE_PHC4060_n2221 (.Y(FE_PHN4060_n2221), 
	.A(n2221));
   DLY4X1 FE_PHC4059_n1941 (.Y(FE_PHN4059_n1941), 
	.A(n1941));
   DLY4X1 FE_PHC4058_n1395 (.Y(FE_PHN4058_n1395), 
	.A(n1395));
   DLY4X1 FE_PHC4057_n991 (.Y(FE_PHN4057_n991), 
	.A(n991));
   DLY4X1 FE_PHC4056_n1519 (.Y(FE_PHN4056_n1519), 
	.A(n1519));
   DLY4X1 FE_PHC4055_n1725 (.Y(FE_PHN4055_n1725), 
	.A(n1725));
   DLY4X1 FE_PHC4054_n2279 (.Y(FE_PHN4054_n2279), 
	.A(n2279));
   DLY4X1 FE_PHC4053_n2000 (.Y(FE_PHN4053_n2000), 
	.A(n2000));
   DLY4X1 FE_PHC4052_n1055 (.Y(FE_PHN4052_n1055), 
	.A(n1055));
   DLY4X1 FE_PHC4051_n2122 (.Y(FE_PHN4051_n2122), 
	.A(n2122));
   DLY4X1 FE_PHC4050_n2085 (.Y(FE_PHN4050_n2085), 
	.A(n2085));
   DLY4X1 FE_PHC4049_n2063 (.Y(FE_PHN4049_n2063), 
	.A(n2063));
   DLY4X1 FE_PHC4048_n890 (.Y(FE_PHN4048_n890), 
	.A(n890));
   DLY4X1 FE_PHC4047_n1185 (.Y(FE_PHN4047_n1185), 
	.A(n1185));
   DLY4X1 FE_PHC4046_n966 (.Y(FE_PHN4046_n966), 
	.A(n966));
   DLY4X1 FE_PHC4045_n1578 (.Y(FE_PHN4045_n1578), 
	.A(n1578));
   DLY4X1 FE_PHC4044_n1646 (.Y(FE_PHN4044_n1646), 
	.A(n1646));
   DLY4X1 FE_PHC4043_n1740 (.Y(FE_PHN4043_n1740), 
	.A(n1740));
   DLY4X1 FE_PHC4042_n1928 (.Y(FE_PHN4042_n1928), 
	.A(n1928));
   DLY4X1 FE_PHC4041_n996 (.Y(FE_PHN4041_n996), 
	.A(n996));
   DLY4X1 FE_PHC4040_n1023 (.Y(FE_PHN4040_n1023), 
	.A(n1023));
   DLY4X1 FE_PHC4039_n950 (.Y(FE_PHN4039_n950), 
	.A(n950));
   DLY4X1 FE_PHC4038_n1515 (.Y(FE_PHN4038_n1515), 
	.A(n1515));
   DLY4X1 FE_PHC4037_n1466 (.Y(FE_PHN4037_n1466), 
	.A(n1466));
   DLY4X1 FE_PHC4036_n1866 (.Y(FE_PHN4036_n1866), 
	.A(n1866));
   DLY4X1 FE_PHC4035_n1544 (.Y(FE_PHN4035_n1544), 
	.A(n1544));
   DLY4X1 FE_PHC4034_n2285 (.Y(FE_PHN4034_n2285), 
	.A(n2285));
   DLY4X1 FE_PHC4033_n2101 (.Y(FE_PHN4033_n2101), 
	.A(n2101));
   DLY4X1 FE_PHC4032_n1012 (.Y(FE_PHN4032_n1012), 
	.A(n1012));
   DLY4X1 FE_PHC4031_n1403 (.Y(FE_PHN4031_n1403), 
	.A(n1403));
   DLY4X1 FE_PHC4030_n1757 (.Y(FE_PHN4030_n1757), 
	.A(n1757));
   DLY4X1 FE_PHC4029_n2100 (.Y(FE_PHN4029_n2100), 
	.A(n2100));
   DLY4X1 FE_PHC4028_n2028 (.Y(FE_PHN4028_n2028), 
	.A(n2028));
   DLY4X1 FE_PHC4027_n2386 (.Y(FE_PHN4027_n2386), 
	.A(n2386));
   DLY4X1 FE_PHC4026_n1741 (.Y(FE_PHN4026_n1741), 
	.A(n1741));
   DLY4X1 FE_PHC4025_n1128 (.Y(FE_PHN4025_n1128), 
	.A(n1128));
   DLY4X1 FE_PHC4024_n986 (.Y(FE_PHN4024_n986), 
	.A(n986));
   DLY4X1 FE_PHC4023_n1854 (.Y(FE_PHN4023_n1854), 
	.A(n1854));
   DLY4X1 FE_PHC4022_n2281 (.Y(FE_PHN4022_n2281), 
	.A(n2281));
   DLY4X1 FE_PHC4021_n2237 (.Y(FE_PHN4021_n2237), 
	.A(n2237));
   DLY4X1 FE_PHC4020_n1547 (.Y(FE_PHN4020_n1547), 
	.A(n1547));
   DLY4X1 FE_PHC4019_n1314 (.Y(FE_PHN4019_n1314), 
	.A(n1314));
   DLY4X1 FE_PHC4018_n944 (.Y(FE_PHN4018_n944), 
	.A(n944));
   DLY4X1 FE_PHC4017_n1456 (.Y(FE_PHN4017_n1456), 
	.A(n1456));
   DLY4X1 FE_PHC4016_n1919 (.Y(FE_PHN4016_n1919), 
	.A(n1919));
   DLY4X1 FE_PHC4015_n897 (.Y(FE_PHN4015_n897), 
	.A(n897));
   DLY4X1 FE_PHC4014_n1297 (.Y(FE_PHN4014_n1297), 
	.A(n1297));
   DLY4X1 FE_PHC4013_n1495 (.Y(FE_PHN4013_n1495), 
	.A(n1495));
   DLY4X1 FE_PHC4012_n1600 (.Y(FE_PHN4012_n1600), 
	.A(n1600));
   DLY4X1 FE_PHC4011_n2102 (.Y(FE_PHN4011_n2102), 
	.A(n2102));
   DLY4X1 FE_PHC4010_n1143 (.Y(FE_PHN4010_n1143), 
	.A(n1143));
   DLY4X1 FE_PHC4009_n2135 (.Y(FE_PHN4009_n2135), 
	.A(n2135));
   DLY4X1 FE_PHC4008_n1474 (.Y(FE_PHN4008_n1474), 
	.A(n1474));
   DLY4X1 FE_PHC4007_n1704 (.Y(FE_PHN4007_n1704), 
	.A(n1704));
   DLY4X1 FE_PHC4006_n1522 (.Y(FE_PHN4006_n1522), 
	.A(n1522));
   DLY4X1 FE_PHC4005_n2162 (.Y(FE_PHN4005_n2162), 
	.A(n2162));
   DLY4X1 FE_PHC4004_n2048 (.Y(FE_PHN4004_n2048), 
	.A(n2048));
   DLY4X1 FE_PHC4003_n894 (.Y(FE_PHN4003_n894), 
	.A(n894));
   DLY4X1 FE_PHC4002_n1382 (.Y(FE_PHN4002_n1382), 
	.A(n1382));
   DLY4X1 FE_PHC4001_n949 (.Y(FE_PHN4001_n949), 
	.A(n949));
   DLY4X1 FE_PHC4000_n1875 (.Y(FE_PHN4000_n1875), 
	.A(n1875));
   DLY4X1 FE_PHC3999_n1896 (.Y(FE_PHN3999_n1896), 
	.A(n1896));
   DLY4X1 FE_PHC3998_n1890 (.Y(FE_PHN3998_n1890), 
	.A(n1890));
   DLY4X1 FE_PHC3997_n2252 (.Y(FE_PHN3997_n2252), 
	.A(n2252));
   DLY4X1 FE_PHC3996_n2096 (.Y(FE_PHN3996_n2096), 
	.A(n2096));
   DLY4X1 FE_PHC3995_n2257 (.Y(FE_PHN3995_n2257), 
	.A(n2257));
   DLY4X1 FE_PHC3994_n1310 (.Y(FE_PHN3994_n1310), 
	.A(n1310));
   DLY4X1 FE_PHC3993_n1367 (.Y(FE_PHN3993_n1367), 
	.A(n1367));
   DLY4X1 FE_PHC3992_n1175 (.Y(FE_PHN3992_n1175), 
	.A(n1175));
   DLY4X1 FE_PHC3991_n2066 (.Y(FE_PHN3991_n2066), 
	.A(n2066));
   DLY4X1 FE_PHC3990_n2268 (.Y(FE_PHN3990_n2268), 
	.A(n2268));
   DLY4X1 FE_PHC3989_n1467 (.Y(FE_PHN3989_n1467), 
	.A(n1467));
   DLY4X1 FE_PHC3988_n2262 (.Y(FE_PHN3988_n2262), 
	.A(n2262));
   DLY3X1 FE_PHC3987_n1686 (.Y(FE_PHN3987_n1686), 
	.A(n1686));
   DLY4X1 FE_PHC3986_n946 (.Y(FE_PHN3986_n946), 
	.A(n946));
   DLY4X1 FE_PHC3985_n2127 (.Y(FE_PHN3985_n2127), 
	.A(n2127));
   DLY4X1 FE_PHC3984_n1483 (.Y(FE_PHN3984_n1483), 
	.A(n1483));
   DLY4X1 FE_PHC3983_n1844 (.Y(FE_PHN3983_n1844), 
	.A(n1844));
   DLY4X1 FE_PHC3982_n2095 (.Y(FE_PHN3982_n2095), 
	.A(n2095));
   DLY4X1 FE_PHC3981_n1850 (.Y(FE_PHN3981_n1850), 
	.A(n1850));
   DLY4X1 FE_PHC3980_n1957 (.Y(FE_PHN3980_n1957), 
	.A(n1957));
   DLY4X1 FE_PHC3979_n1948 (.Y(FE_PHN3979_n1948), 
	.A(n1948));
   DLY4X1 FE_PHC3978_n972 (.Y(FE_PHN3978_n972), 
	.A(n972));
   DLY4X1 FE_PHC3977_n903 (.Y(FE_PHN3977_n903), 
	.A(n903));
   DLY4X1 FE_PHC3976_n982 (.Y(FE_PHN3976_n982), 
	.A(n982));
   DLY4X1 FE_PHC3975_n1400 (.Y(FE_PHN3975_n1400), 
	.A(n1400));
   DLY4X1 FE_PHC3974_n1846 (.Y(FE_PHN3974_n1846), 
	.A(n1846));
   DLY4X1 FE_PHC3973_n1402 (.Y(FE_PHN3973_n1402), 
	.A(n1402));
   DLY4X1 FE_PHC3972_n2110 (.Y(FE_PHN3972_n2110), 
	.A(n2110));
   DLY4X1 FE_PHC3971_n1698 (.Y(FE_PHN3971_n1698), 
	.A(n1698));
   DLY4X1 FE_PHC3970_n1680 (.Y(FE_PHN3970_n1680), 
	.A(n1680));
   DLY4X1 FE_PHC3969_n1696 (.Y(FE_PHN3969_n1696), 
	.A(n1696));
   DLY4X1 FE_PHC3968_n1664 (.Y(FE_PHN3968_n1664), 
	.A(n1664));
   DLY4X1 FE_PHC3967_n1114 (.Y(FE_PHN3967_n1114), 
	.A(n1114));
   DLY4X1 FE_PHC3966_n1433 (.Y(FE_PHN3966_n1433), 
	.A(n1433));
   DLY4X1 FE_PHC3965_n1476 (.Y(FE_PHN3965_n1476), 
	.A(n1476));
   DLY4X1 FE_PHC3964_n1715 (.Y(FE_PHN3964_n1715), 
	.A(n1715));
   DLY4X1 FE_PHC3963_n905 (.Y(FE_PHN3963_n905), 
	.A(n905));
   DLY4X1 FE_PHC3962_n1772 (.Y(FE_PHN3962_n1772), 
	.A(n1772));
   DLY4X1 FE_PHC3961_n2006 (.Y(FE_PHN3961_n2006), 
	.A(n2006));
   DLY4X1 FE_PHC3960_n1549 (.Y(FE_PHN3960_n1549), 
	.A(n1549));
   DLY4X1 FE_PHC3959_n2108 (.Y(FE_PHN3959_n2108), 
	.A(n2108));
   DLY4X1 FE_PHC3958_n2034 (.Y(FE_PHN3958_n2034), 
	.A(n2034));
   DLY4X1 FE_PHC3957_n951 (.Y(FE_PHN3957_n951), 
	.A(n951));
   DLY4X1 FE_PHC3956_n955 (.Y(FE_PHN3956_n955), 
	.A(n955));
   DLY4X1 FE_PHC3955_n1709 (.Y(FE_PHN3955_n1709), 
	.A(n1709));
   DLY4X1 FE_PHC3954_n2183 (.Y(FE_PHN3954_n2183), 
	.A(n2183));
   DLY4X1 FE_PHC3953_n2211 (.Y(FE_PHN3953_n2211), 
	.A(n2211));
   DLY4X1 FE_PHC3952_n1868 (.Y(FE_PHN3952_n1868), 
	.A(n1868));
   DLY4X1 FE_PHC3951_n1913 (.Y(FE_PHN3951_n1913), 
	.A(n1913));
   DLY4X1 FE_PHC3950_n1521 (.Y(FE_PHN3950_n1521), 
	.A(n1521));
   DLY4X1 FE_PHC3949_n1576 (.Y(FE_PHN3949_n1576), 
	.A(n1576));
   DLY4X1 FE_PHC3948_n1789 (.Y(FE_PHN3948_n1789), 
	.A(n1789));
   DLY4X1 FE_PHC3947_n1316 (.Y(FE_PHN3947_n1316), 
	.A(n1316));
   DLY4X1 FE_PHC3946_n1815 (.Y(FE_PHN3946_n1815), 
	.A(n1815));
   DLY4X1 FE_PHC3945_n1821 (.Y(FE_PHN3945_n1821), 
	.A(n1821));
   DLY4X1 FE_PHC3944_n2192 (.Y(FE_PHN3944_n2192), 
	.A(n2192));
   DLY4X1 FE_PHC3943_n2272 (.Y(FE_PHN3943_n2272), 
	.A(n2272));
   DLY4X1 FE_PHC3942_n922 (.Y(FE_PHN3942_n922), 
	.A(n922));
   DLY4X1 FE_PHC3941_n985 (.Y(FE_PHN3941_n985), 
	.A(n985));
   DLY4X1 FE_PHC3940_n1795 (.Y(FE_PHN3940_n1795), 
	.A(n1795));
   DLY4X1 FE_PHC3939_n1000 (.Y(FE_PHN3939_n1000), 
	.A(n1000));
   DLY4X1 FE_PHC3938_n1824 (.Y(FE_PHN3938_n1824), 
	.A(n1824));
   DLY4X1 FE_PHC3937_n1747 (.Y(FE_PHN3937_n1747), 
	.A(n1747));
   DLY4X1 FE_PHC3936_n2246 (.Y(FE_PHN3936_n2246), 
	.A(n2246));
   DLY4X1 FE_PHC3935_n2109 (.Y(FE_PHN3935_n2109), 
	.A(n2109));
   DLY4X1 FE_PHC3934_n1739 (.Y(FE_PHN3934_n1739), 
	.A(n1739));
   DLY4X1 FE_PHC3933_n1580 (.Y(FE_PHN3933_n1580), 
	.A(n1580));
   DLY4X1 FE_PHC3932_n1804 (.Y(FE_PHN3932_n1804), 
	.A(n1804));
   DLY4X1 FE_PHC3931_n2249 (.Y(FE_PHN3931_n2249), 
	.A(n2249));
   DLY4X1 FE_PHC3930_n2142 (.Y(FE_PHN3930_n2142), 
	.A(n2142));
   DLY4X1 FE_PHC3929_n1802 (.Y(FE_PHN3929_n1802), 
	.A(n1802));
   DLY4X1 FE_PHC3928_n1041 (.Y(FE_PHN3928_n1041), 
	.A(n1041));
   DLY4X1 FE_PHC3927_n930 (.Y(FE_PHN3927_n930), 
	.A(n930));
   DLY4X1 FE_PHC3926_n1869 (.Y(FE_PHN3926_n1869), 
	.A(n1869));
   DLY4X1 FE_PHC3925_n1699 (.Y(FE_PHN3925_n1699), 
	.A(n1699));
   DLY4X1 FE_PHC3924_n1524 (.Y(FE_PHN3924_n1524), 
	.A(n1524));
   DLY4X1 FE_PHC3923_n2087 (.Y(FE_PHN3923_n2087), 
	.A(n2087));
   DLY4X1 FE_PHC3922_n1397 (.Y(FE_PHN3922_n1397), 
	.A(n1397));
   DLY4X1 FE_PHC3921_n1459 (.Y(FE_PHN3921_n1459), 
	.A(n1459));
   DLY4X1 FE_PHC3920_n1441 (.Y(FE_PHN3920_n1441), 
	.A(n1441));
   DLY4X1 FE_PHC3919_n967 (.Y(FE_PHN3919_n967), 
	.A(n967));
   DLY4X1 FE_PHC3918_n1684 (.Y(FE_PHN3918_n1684), 
	.A(n1684));
   DLY4X1 FE_PHC3917_n1921 (.Y(FE_PHN3917_n1921), 
	.A(n1921));
   DLY4X1 FE_PHC3916_n2062 (.Y(FE_PHN3916_n2062), 
	.A(n2062));
   DLY3X1 FE_PHC3915_n2168 (.Y(FE_PHN3915_n2168), 
	.A(n2168));
   DLY4X1 FE_PHC3914_n2041 (.Y(FE_PHN3914_n2041), 
	.A(n2041));
   DLY4X1 FE_PHC3913_n1858 (.Y(FE_PHN3913_n1858), 
	.A(n1858));
   DLY4X1 FE_PHC3912_n1876 (.Y(FE_PHN3912_n1876), 
	.A(n1876));
   DLY4X1 FE_PHC3911_n1428 (.Y(FE_PHN3911_n1428), 
	.A(n1428));
   DLY4X1 FE_PHC3910_n1431 (.Y(FE_PHN3910_n1431), 
	.A(n1431));
   DLY4X1 FE_PHC3909_n2001 (.Y(FE_PHN3909_n2001), 
	.A(n2001));
   DLY4X1 FE_PHC3908_n2243 (.Y(FE_PHN3908_n2243), 
	.A(n2243));
   DLY4X1 FE_PHC3907_n1491 (.Y(FE_PHN3907_n1491), 
	.A(n1491));
   DLY4X1 FE_PHC3906_n1877 (.Y(FE_PHN3906_n1877), 
	.A(n1877));
   DLY4X1 FE_PHC3905_n1883 (.Y(FE_PHN3905_n1883), 
	.A(n1883));
   DLY4X1 FE_PHC3904_n1702 (.Y(FE_PHN3904_n1702), 
	.A(n1702));
   DLY4X1 FE_PHC3903_n2143 (.Y(FE_PHN3903_n2143), 
	.A(n2143));
   DLY4X1 FE_PHC3902_n1703 (.Y(FE_PHN3902_n1703), 
	.A(n1703));
   DLY4X1 FE_PHC3901_n1711 (.Y(FE_PHN3901_n1711), 
	.A(n1711));
   DLY4X1 FE_PHC3900_n2082 (.Y(FE_PHN3900_n2082), 
	.A(n2082));
   DLY4X1 FE_PHC3899_n2118 (.Y(FE_PHN3899_n2118), 
	.A(n2118));
   DLY4X1 FE_PHC3898_n2170 (.Y(FE_PHN3898_n2170), 
	.A(n2170));
   DLY4X1 FE_PHC3897_n1448 (.Y(FE_PHN3897_n1448), 
	.A(n1448));
   DLY4X1 FE_PHC3896_n1797 (.Y(FE_PHN3896_n1797), 
	.A(n1797));
   DLY4X1 FE_PHC3895_n2051 (.Y(FE_PHN3895_n2051), 
	.A(n2051));
   DLY4X1 FE_PHC3894_n1874 (.Y(FE_PHN3894_n1874), 
	.A(n1874));
   DLY4X1 FE_PHC3893_n2286 (.Y(FE_PHN3893_n2286), 
	.A(n2286));
   DLY4X1 FE_PHC3892_n1759 (.Y(FE_PHN3892_n1759), 
	.A(n1759));
   DLY4X1 FE_PHC3891_n2072 (.Y(FE_PHN3891_n2072), 
	.A(n2072));
   DLY4X1 FE_PHC3890_n1807 (.Y(FE_PHN3890_n1807), 
	.A(n1807));
   DLY4X1 FE_PHC3889_n2077 (.Y(FE_PHN3889_n2077), 
	.A(n2077));
   DLY4X1 FE_PHC3888_n2254 (.Y(FE_PHN3888_n2254), 
	.A(n2254));
   DLY4X1 FE_PHC3887_n1701 (.Y(FE_PHN3887_n1701), 
	.A(n1701));
   DLY4X1 FE_PHC3886_n2103 (.Y(FE_PHN3886_n2103), 
	.A(n2103));
   DLY4X1 FE_PHC3885_n1768 (.Y(FE_PHN3885_n1768), 
	.A(n1768));
   DLY4X1 FE_PHC3884_n923 (.Y(FE_PHN3884_n923), 
	.A(n923));
   DLY4X1 FE_PHC3883_n1594 (.Y(FE_PHN3883_n1594), 
	.A(n1594));
   DLY4X1 FE_PHC3882_n2230 (.Y(FE_PHN3882_n2230), 
	.A(n2230));
   DLY4X1 FE_PHC3881_n1481 (.Y(FE_PHN3881_n1481), 
	.A(n1481));
   DLY4X1 FE_PHC3880_n938 (.Y(FE_PHN3880_n938), 
	.A(n938));
   DLY4X1 FE_PHC3879_n1497 (.Y(FE_PHN3879_n1497), 
	.A(n1497));
   DLY4X1 FE_PHC3878_n1852 (.Y(FE_PHN3878_n1852), 
	.A(n1852));
   DLY4X1 FE_PHC3877_n889 (.Y(FE_PHN3877_n889), 
	.A(n889));
   DLY4X1 FE_PHC3876_n2205 (.Y(FE_PHN3876_n2205), 
	.A(n2205));
   DLY4X1 FE_PHC3875_n1829 (.Y(FE_PHN3875_n1829), 
	.A(n1829));
   DLY4X1 FE_PHC3874_n2244 (.Y(FE_PHN3874_n2244), 
	.A(n2244));
   DLY4X1 FE_PHC3873_n2270 (.Y(FE_PHN3873_n2270), 
	.A(n2270));
   DLY4X1 FE_PHC3872_n1778 (.Y(FE_PHN3872_n1778), 
	.A(n1778));
   DLY4X1 FE_PHC3871_n1655 (.Y(FE_PHN3871_n1655), 
	.A(n1655));
   DLY4X1 FE_PHC3870_n2208 (.Y(FE_PHN3870_n2208), 
	.A(n2208));
   DLY4X1 FE_PHC3869_n962 (.Y(FE_PHN3869_n962), 
	.A(n962));
   DLY4X1 FE_PHC3868_n1472 (.Y(FE_PHN3868_n1472), 
	.A(n1472));
   DLY4X1 FE_PHC3867_n1762 (.Y(FE_PHN3867_n1762), 
	.A(n1762));
   DLY4X1 FE_PHC3866_n908 (.Y(FE_PHN3866_n908), 
	.A(n908));
   DLY4X1 FE_PHC3865_n1786 (.Y(FE_PHN3865_n1786), 
	.A(n1786));
   DLY4X1 FE_PHC3864_n1738 (.Y(FE_PHN3864_n1738), 
	.A(n1738));
   DLY4X1 FE_PHC3863_n2088 (.Y(FE_PHN3863_n2088), 
	.A(n2088));
   DLY4X1 FE_PHC3862_n1743 (.Y(FE_PHN3862_n1743), 
	.A(n1743));
   DLY4X1 FE_PHC3861_n2068 (.Y(FE_PHN3861_n2068), 
	.A(n2068));
   DLY4X1 FE_PHC3860_n2173 (.Y(FE_PHN3860_n2173), 
	.A(n2173));
   DLY4X1 FE_PHC3859_n1506 (.Y(FE_PHN3859_n1506), 
	.A(n1506));
   DLY4X1 FE_PHC3858_n2374 (.Y(FE_PHN3858_n2374), 
	.A(n2374));
   DLY4X1 FE_PHC3857_n1714 (.Y(FE_PHN3857_n1714), 
	.A(n1714));
   DLY4X1 FE_PHC3856_n1998 (.Y(FE_PHN3856_n1998), 
	.A(n1998));
   DLY4X1 FE_PHC3855_n1631 (.Y(FE_PHN3855_n1631), 
	.A(n1631));
   DLY4X1 FE_PHC3854_n1710 (.Y(FE_PHN3854_n1710), 
	.A(n1710));
   DLY4X1 FE_PHC3853_n964 (.Y(FE_PHN3853_n964), 
	.A(n964));
   DLY4X1 FE_PHC3852_n2225 (.Y(FE_PHN3852_n2225), 
	.A(n2225));
   DLY4X1 FE_PHC3851_n1691 (.Y(FE_PHN3851_n1691), 
	.A(n1691));
   DLY4X1 FE_PHC3850_n1369 (.Y(FE_PHN3850_n1369), 
	.A(n1369));
   DLY4X1 FE_PHC3849_n2245 (.Y(FE_PHN3849_n2245), 
	.A(n2245));
   DLY4X1 FE_PHC3848_n2169 (.Y(FE_PHN3848_n2169), 
	.A(n2169));
   DLY4X1 FE_PHC3847_n2199 (.Y(FE_PHN3847_n2199), 
	.A(n2199));
   DLY4X1 FE_PHC3846_n1939 (.Y(FE_PHN3846_n1939), 
	.A(n1939));
   DLY4X1 FE_PHC3845_n980 (.Y(FE_PHN3845_n980), 
	.A(n980));
   DLY4X1 FE_PHC3844_n1498 (.Y(FE_PHN3844_n1498), 
	.A(n1498));
   DLY4X1 FE_PHC3843_n2233 (.Y(FE_PHN3843_n2233), 
	.A(n2233));
   DLY4X1 FE_PHC3842_n1499 (.Y(FE_PHN3842_n1499), 
	.A(n1499));
   DLY4X1 FE_PHC3841_n1855 (.Y(FE_PHN3841_n1855), 
	.A(n1855));
   DLY4X1 FE_PHC3840_n1523 (.Y(FE_PHN3840_n1523), 
	.A(n1523));
   DLY4X1 FE_PHC3839_n1842 (.Y(FE_PHN3839_n1842), 
	.A(n1842));
   DLY4X1 FE_PHC3838_n1417 (.Y(FE_PHN3838_n1417), 
	.A(n1417));
   DLY4X1 FE_PHC3837_n1873 (.Y(FE_PHN3837_n1873), 
	.A(n1873));
   DLY4X1 FE_PHC3836_n2132 (.Y(FE_PHN3836_n2132), 
	.A(n2132));
   DLY4X1 FE_PHC3835_n1489 (.Y(FE_PHN3835_n1489), 
	.A(n1489));
   DLY4X1 FE_PHC3834_n1490 (.Y(FE_PHN3834_n1490), 
	.A(n1490));
   DLY4X1 FE_PHC3833_n1437 (.Y(FE_PHN3833_n1437), 
	.A(n1437));
   DLY4X1 FE_PHC3832_n2075 (.Y(FE_PHN3832_n2075), 
	.A(n2075));
   DLY4X1 FE_PHC3831_n2177 (.Y(FE_PHN3831_n2177), 
	.A(n2177));
   DLY4X1 FE_PHC3830_n1593 (.Y(FE_PHN3830_n1593), 
	.A(n1593));
   DLY4X1 FE_PHC3829_n1577 (.Y(FE_PHN3829_n1577), 
	.A(n1577));
   DLY4X1 FE_PHC3828_n2203 (.Y(FE_PHN3828_n2203), 
	.A(n2203));
   DLY4X1 FE_PHC3827_n1492 (.Y(FE_PHN3827_n1492), 
	.A(n1492));
   DLY4X1 FE_PHC3826_n1870 (.Y(FE_PHN3826_n1870), 
	.A(n1870));
   DLY4X1 FE_PHC3825_n1618 (.Y(FE_PHN3825_n1618), 
	.A(n1618));
   DLY4X1 FE_PHC3824_n1835 (.Y(FE_PHN3824_n1835), 
	.A(n1835));
   DLY4X1 FE_PHC3823_n2067 (.Y(FE_PHN3823_n2067), 
	.A(n2067));
   DLY4X1 FE_PHC3822_n1894 (.Y(FE_PHN3822_n1894), 
	.A(n1894));
   DLY4X1 FE_PHC3821_n1555 (.Y(FE_PHN3821_n1555), 
	.A(n1555));
   DLY4X1 FE_PHC3820_n1415 (.Y(FE_PHN3820_n1415), 
	.A(n1415));
   DLY4X1 FE_PHC3819_n2372 (.Y(FE_PHN3819_n2372), 
	.A(n2372));
   DLY4X1 FE_PHC3818_n898 (.Y(FE_PHN3818_n898), 
	.A(n898));
   DLY4X1 FE_PHC3817_n1745 (.Y(FE_PHN3817_n1745), 
	.A(n1745));
   DLY4X1 FE_PHC3816_n1662 (.Y(FE_PHN3816_n1662), 
	.A(n1662));
   DLY4X1 FE_PHC3815_n1880 (.Y(FE_PHN3815_n1880), 
	.A(n1880));
   DLY4X1 FE_PHC3814_n2210 (.Y(FE_PHN3814_n2210), 
	.A(n2210));
   DLY4X1 FE_PHC3813_n1672 (.Y(FE_PHN3813_n1672), 
	.A(n1672));
   DLY4X1 FE_PHC3812_n1822 (.Y(FE_PHN3812_n1822), 
	.A(n1822));
   DLY4X1 FE_PHC3811_n2265 (.Y(FE_PHN3811_n2265), 
	.A(n2265));
   DLY4X1 FE_PHC3810_n1906 (.Y(FE_PHN3810_n1906), 
	.A(n1906));
   DLY4X1 FE_PHC3809_n2269 (.Y(FE_PHN3809_n2269), 
	.A(n2269));
   DLY4X1 FE_PHC3808_n1781 (.Y(FE_PHN3808_n1781), 
	.A(n1781));
   DLY4X1 FE_PHC3807_n2214 (.Y(FE_PHN3807_n2214), 
	.A(n2214));
   DLY4X1 FE_PHC3806_n2130 (.Y(FE_PHN3806_n2130), 
	.A(n2130));
   DLY4X1 FE_PHC3805_n1673 (.Y(FE_PHN3805_n1673), 
	.A(n1673));
   DLY4X1 FE_PHC3804_n2080 (.Y(FE_PHN3804_n2080), 
	.A(n2080));
   DLY4X1 FE_PHC3803_n1473 (.Y(FE_PHN3803_n1473), 
	.A(n1473));
   DLY4X1 FE_PHC3802_n2150 (.Y(FE_PHN3802_n2150), 
	.A(n2150));
   DLY4X1 FE_PHC3801_n1502 (.Y(FE_PHN3801_n1502), 
	.A(n1502));
   DLY4X1 FE_PHC3800_n1898 (.Y(FE_PHN3800_n1898), 
	.A(n1898));
   DLY4X1 FE_PHC3799_n1723 (.Y(FE_PHN3799_n1723), 
	.A(n1723));
   DLY4X1 FE_PHC3798_n1597 (.Y(FE_PHN3798_n1597), 
	.A(n1597));
   DLY4X1 FE_PHC3797_n893 (.Y(FE_PHN3797_n893), 
	.A(n893));
   DLY4X1 FE_PHC3796_n2086 (.Y(FE_PHN3796_n2086), 
	.A(n2086));
   DLY4X1 FE_PHC3795_n1486 (.Y(FE_PHN3795_n1486), 
	.A(n1486));
   DLY4X1 FE_PHC3794_n1604 (.Y(FE_PHN3794_n1604), 
	.A(n1604));
   DLY4X1 FE_PHC3793_n1719 (.Y(FE_PHN3793_n1719), 
	.A(n1719));
   DLY4X1 FE_PHC3792_n1438 (.Y(FE_PHN3792_n1438), 
	.A(n1438));
   DLY4X1 FE_PHC3791_n2089 (.Y(FE_PHN3791_n2089), 
	.A(n2089));
   DLY4X1 FE_PHC3790_n1817 (.Y(FE_PHN3790_n1817), 
	.A(n1817));
   DLY4X1 FE_PHC3789_n1750 (.Y(FE_PHN3789_n1750), 
	.A(n1750));
   DLY4X1 FE_PHC3788_n1399 (.Y(FE_PHN3788_n1399), 
	.A(n1399));
   DLY4X1 FE_PHC3787_n1805 (.Y(FE_PHN3787_n1805), 
	.A(n1805));
   DLY4X1 FE_PHC3786_n1945 (.Y(FE_PHN3786_n1945), 
	.A(n1945));
   DLY4X1 FE_PHC3785_n2276 (.Y(FE_PHN3785_n2276), 
	.A(n2276));
   DLY4X1 FE_PHC3784_n1657 (.Y(FE_PHN3784_n1657), 
	.A(n1657));
   DLY4X1 FE_PHC3783_n2202 (.Y(FE_PHN3783_n2202), 
	.A(n2202));
   DLY4X1 FE_PHC3782_n1364 (.Y(FE_PHN3782_n1364), 
	.A(n1364));
   DLY4X1 FE_PHC3781_n1727 (.Y(FE_PHN3781_n1727), 
	.A(n1727));
   DLY4X1 FE_PHC3780_n2213 (.Y(FE_PHN3780_n2213), 
	.A(n2213));
   DLY4X1 FE_PHC3779_n1726 (.Y(FE_PHN3779_n1726), 
	.A(n1726));
   DLY4X1 FE_PHC3778_n2079 (.Y(FE_PHN3778_n2079), 
	.A(n2079));
   DLY4X1 FE_PHC3777_n2097 (.Y(FE_PHN3777_n2097), 
	.A(n2097));
   DLY4X1 FE_PHC3776_n1660 (.Y(FE_PHN3776_n1660), 
	.A(n1660));
   DLY4X1 FE_PHC3775_n1509 (.Y(FE_PHN3775_n1509), 
	.A(n1509));
   DLY4X1 FE_PHC3774_n1967 (.Y(FE_PHN3774_n1967), 
	.A(n1967));
   DLY4X1 FE_PHC3773_n1404 (.Y(FE_PHN3773_n1404), 
	.A(n1404));
   DLY4X1 FE_PHC3772_n1756 (.Y(FE_PHN3772_n1756), 
	.A(n1756));
   DLY4X1 FE_PHC3771_n1508 (.Y(FE_PHN3771_n1508), 
	.A(n1508));
   DLY4X1 FE_PHC3770_n1860 (.Y(FE_PHN3770_n1860), 
	.A(n1860));
   DLY4X1 FE_PHC3769_n1705 (.Y(FE_PHN3769_n1705), 
	.A(n1705));
   DLY4X1 FE_PHC3768_n1729 (.Y(FE_PHN3768_n1729), 
	.A(n1729));
   DLY4X1 FE_PHC3767_n1465 (.Y(FE_PHN3767_n1465), 
	.A(n1465));
   DLY4X1 FE_PHC3766_n1882 (.Y(FE_PHN3766_n1882), 
	.A(n1882));
   DLY4X1 FE_PHC3765_n2259 (.Y(FE_PHN3765_n2259), 
	.A(n2259));
   DLY4X1 FE_PHC3764_n2083 (.Y(FE_PHN3764_n2083), 
	.A(n2083));
   DLY4X1 FE_PHC3763_n2044 (.Y(FE_PHN3763_n2044), 
	.A(n2044));
   DLY4X1 FE_PHC3762_n2055 (.Y(FE_PHN3762_n2055), 
	.A(n2055));
   DLY4X1 FE_PHC3761_n1760 (.Y(FE_PHN3761_n1760), 
	.A(n1760));
   DLY4X1 FE_PHC3760_n1671 (.Y(FE_PHN3760_n1671), 
	.A(n1671));
   DLY4X1 FE_PHC3759_n1494 (.Y(FE_PHN3759_n1494), 
	.A(n1494));
   DLY4X1 FE_PHC3758_n1871 (.Y(FE_PHN3758_n1871), 
	.A(n1871));
   DLY4X1 FE_PHC3757_n1754 (.Y(FE_PHN3757_n1754), 
	.A(n1754));
   DLY4X1 FE_PHC3756_n1443 (.Y(FE_PHN3756_n1443), 
	.A(n1443));
   DLY4X1 FE_PHC3755_n1769 (.Y(FE_PHN3755_n1769), 
	.A(n1769));
   DLY4X1 FE_PHC3754_n2198 (.Y(FE_PHN3754_n2198), 
	.A(n2198));
   DLY4X1 FE_PHC3753_n1406 (.Y(FE_PHN3753_n1406), 
	.A(n1406));
   DLY4X1 FE_PHC3752_n1798 (.Y(FE_PHN3752_n1798), 
	.A(n1798));
   DLY4X1 FE_PHC3751_n2227 (.Y(FE_PHN3751_n2227), 
	.A(n2227));
   DLY4X1 FE_PHC3750_n1801 (.Y(FE_PHN3750_n1801), 
	.A(n1801));
   DLY4X1 FE_PHC3749_n1458 (.Y(FE_PHN3749_n1458), 
	.A(n1458));
   DLY4X1 FE_PHC3748_n1787 (.Y(FE_PHN3748_n1787), 
	.A(n1787));
   DLY4X1 FE_PHC3747_n1411 (.Y(FE_PHN3747_n1411), 
	.A(n1411));
   DLY4X1 FE_PHC3746_n2178 (.Y(FE_PHN3746_n2178), 
	.A(n2178));
   DLY4X1 FE_PHC3745_n2078 (.Y(FE_PHN3745_n2078), 
	.A(n2078));
   DLY4X1 FE_PHC3744_n1803 (.Y(FE_PHN3744_n1803), 
	.A(n1803));
   DLY4X1 FE_PHC3743_n2069 (.Y(FE_PHN3743_n2069), 
	.A(n2069));
   DLY4X1 FE_PHC3742_n1451 (.Y(FE_PHN3742_n1451), 
	.A(n1451));
   DLY4X1 FE_PHC3741_n2134 (.Y(FE_PHN3741_n2134), 
	.A(n2134));
   DLY4X1 FE_PHC3740_n2242 (.Y(FE_PHN3740_n2242), 
	.A(n2242));
   DLY4X1 FE_PHC3739_n2195 (.Y(FE_PHN3739_n2195), 
	.A(n2195));
   DLY4X1 FE_PHC3738_n1863 (.Y(FE_PHN3738_n1863), 
	.A(n1863));
   DLY4X1 FE_PHC3737_n2098 (.Y(FE_PHN3737_n2098), 
	.A(n2098));
   DLY4X1 FE_PHC3736_n2264 (.Y(FE_PHN3736_n2264), 
	.A(n2264));
   DLY4X1 FE_PHC3735_n1511 (.Y(FE_PHN3735_n1511), 
	.A(n1511));
   DLY4X1 FE_PHC3734_n2054 (.Y(FE_PHN3734_n2054), 
	.A(n2054));
   DLY4X1 FE_PHC3733_n1774 (.Y(FE_PHN3733_n1774), 
	.A(n1774));
   DLY4X1 FE_PHC3732_n2260 (.Y(FE_PHN3732_n2260), 
	.A(n2260));
   DLY4X1 FE_PHC3731_n1444 (.Y(FE_PHN3731_n1444), 
	.A(n1444));
   DLY4X1 FE_PHC3730_n2187 (.Y(FE_PHN3730_n2187), 
	.A(n2187));
   DLY4X1 FE_PHC3729_n2160 (.Y(FE_PHN3729_n2160), 
	.A(n2160));
   DLY4X1 FE_PHC3728_n2251 (.Y(FE_PHN3728_n2251), 
	.A(n2251));
   DLY4X1 FE_PHC3727_n2146 (.Y(FE_PHN3727_n2146), 
	.A(n2146));
   DLY4X1 FE_PHC3726_n1823 (.Y(FE_PHN3726_n1823), 
	.A(n1823));
   DLY4X1 FE_PHC3725_n2145 (.Y(FE_PHN3725_n2145), 
	.A(n2145));
   DLY4X1 FE_PHC3724_n2218 (.Y(FE_PHN3724_n2218), 
	.A(n2218));
   DLY4X1 FE_PHC3723_n1328 (.Y(FE_PHN3723_n1328), 
	.A(n1328));
   DLY4X1 FE_PHC3722_n1840 (.Y(FE_PHN3722_n1840), 
	.A(n1840));
   DLY4X1 FE_PHC3721_n1436 (.Y(FE_PHN3721_n1436), 
	.A(n1436));
   DLY4X1 FE_PHC3720_n1752 (.Y(FE_PHN3720_n1752), 
	.A(n1752));
   DLY4X1 FE_PHC3719_n1721 (.Y(FE_PHN3719_n1721), 
	.A(n1721));
   DLY4X1 FE_PHC3718_n1429 (.Y(FE_PHN3718_n1429), 
	.A(n1429));
   DLY4X1 FE_PHC3717_n2288 (.Y(FE_PHN3717_n2288), 
	.A(n2288));
   DLY4X1 FE_PHC3716_n1439 (.Y(FE_PHN3716_n1439), 
	.A(n1439));
   DLY4X1 FE_PHC3715_n2074 (.Y(FE_PHN3715_n2074), 
	.A(n2074));
   DLY4X1 FE_PHC3714_n2217 (.Y(FE_PHN3714_n2217), 
	.A(n2217));
   DLY4X1 FE_PHC3713_n1424 (.Y(FE_PHN3713_n1424), 
	.A(n1424));
   DLY4X1 FE_PHC3712_n2112 (.Y(FE_PHN3712_n2112), 
	.A(n2112));
   DLY4X1 FE_PHC3711_n2204 (.Y(FE_PHN3711_n2204), 
	.A(n2204));
   DLY4X1 FE_PHC3710_n1656 (.Y(FE_PHN3710_n1656), 
	.A(n1656));
   DLY4X1 FE_PHC3709_n1512 (.Y(FE_PHN3709_n1512), 
	.A(n1512));
   DLY4X1 FE_PHC3708_n2099 (.Y(FE_PHN3708_n2099), 
	.A(n2099));
   DLY4X1 FE_PHC3707_n2129 (.Y(FE_PHN3707_n2129), 
	.A(n2129));
   DLY4X1 FE_PHC3706_n1694 (.Y(FE_PHN3706_n1694), 
	.A(n1694));
   DLY4X1 FE_PHC3705_n2141 (.Y(FE_PHN3705_n2141), 
	.A(n2141));
   DLY4X1 FE_PHC3704_n2224 (.Y(FE_PHN3704_n2224), 
	.A(n2224));
   DLY4X1 FE_PHC3703_n2171 (.Y(FE_PHN3703_n2171), 
	.A(n2171));
   DLY4X1 FE_PHC3702_n2106 (.Y(FE_PHN3702_n2106), 
	.A(n2106));
   DLY4X1 FE_PHC3701_n2175 (.Y(FE_PHN3701_n2175), 
	.A(n2175));
   DLY4X1 FE_PHC3700_n2107 (.Y(FE_PHN3700_n2107), 
	.A(n2107));
   DLY4X1 FE_PHC3699_n1737 (.Y(FE_PHN3699_n1737), 
	.A(n1737));
   DLY4X1 FE_PHC3698_n1722 (.Y(FE_PHN3698_n1722), 
	.A(n1722));
   DLY4X1 FE_PHC3697_n1442 (.Y(FE_PHN3697_n1442), 
	.A(n1442));
   DLY4X1 FE_PHC3696_n1849 (.Y(FE_PHN3696_n1849), 
	.A(n1849));
   DLY4X1 FE_PHC3695_n2250 (.Y(FE_PHN3695_n2250), 
	.A(n2250));
   DLY4X1 FE_PHC3694_n2196 (.Y(FE_PHN3694_n2196), 
	.A(n2196));
   DLY4X1 FE_PHC3693_n2263 (.Y(FE_PHN3693_n2263), 
	.A(n2263));
   DLY4X1 FE_PHC3692_n1667 (.Y(FE_PHN3692_n1667), 
	.A(n1667));
   DLY4X1 FE_PHC3691_n2059 (.Y(FE_PHN3691_n2059), 
	.A(n2059));
   DLY4X1 FE_PHC3690_n1864 (.Y(FE_PHN3690_n1864), 
	.A(n1864));
   DLY4X1 FE_PHC3689_n1904 (.Y(FE_PHN3689_n1904), 
	.A(n1904));
   DLY4X1 FE_PHC3688_n1487 (.Y(FE_PHN3688_n1487), 
	.A(n1487));
   DLY4X1 FE_PHC3687_n1422 (.Y(FE_PHN3687_n1422), 
	.A(n1422));
   DLY4X1 FE_PHC3686_n1814 (.Y(FE_PHN3686_n1814), 
	.A(n1814));
   DLY4X1 FE_PHC3685_n1733 (.Y(FE_PHN3685_n1733), 
	.A(n1733));
   DLY4X1 FE_PHC3684_n1463 (.Y(FE_PHN3684_n1463), 
	.A(n1463));
   DLY4X1 FE_PHC3683_n1893 (.Y(FE_PHN3683_n1893), 
	.A(n1893));
   DLY4X1 FE_PHC3682_n2200 (.Y(FE_PHN3682_n2200), 
	.A(n2200));
   DLY4X1 FE_PHC3681_n1818 (.Y(FE_PHN3681_n1818), 
	.A(n1818));
   DLY4X1 FE_PHC3680_n2206 (.Y(FE_PHN3680_n2206), 
	.A(n2206));
   DLY4X1 FE_PHC3679_n1454 (.Y(FE_PHN3679_n1454), 
	.A(n1454));
   DLY4X1 FE_PHC3678_n2057 (.Y(FE_PHN3678_n2057), 
	.A(n2057));
   DLY4X1 FE_PHC3677_n2190 (.Y(FE_PHN3677_n2190), 
	.A(n2190));
   DLY4X1 FE_PHC3676_n1692 (.Y(FE_PHN3676_n1692), 
	.A(n1692));
   DLY4X1 FE_PHC3675_n1794 (.Y(FE_PHN3675_n1794), 
	.A(n1794));
   DLY4X1 FE_PHC3674_n2092 (.Y(FE_PHN3674_n2092), 
	.A(n2092));
   DLY4X1 FE_PHC3673_n2113 (.Y(FE_PHN3673_n2113), 
	.A(n2113));
   DLY4X1 FE_PHC3672_n2136 (.Y(FE_PHN3672_n2136), 
	.A(n2136));
   DLY4X1 FE_PHC3671_n1687 (.Y(FE_PHN3671_n1687), 
	.A(n1687));
   DLY4X1 FE_PHC3670_n2050 (.Y(FE_PHN3670_n2050), 
	.A(n2050));
   DLY4X1 FE_PHC3669_n1706 (.Y(FE_PHN3669_n1706), 
	.A(n1706));
   DLY4X1 FE_PHC3668_n1452 (.Y(FE_PHN3668_n1452), 
	.A(n1452));
   DLY4X1 FE_PHC3667_n1685 (.Y(FE_PHN3667_n1685), 
	.A(n1685));
   DLY4X1 FE_PHC3666_n1446 (.Y(FE_PHN3666_n1446), 
	.A(n1446));
   DLY4X1 FE_PHC3665_n1764 (.Y(FE_PHN3665_n1764), 
	.A(n1764));
   DLY4X1 FE_PHC3664_n2070 (.Y(FE_PHN3664_n2070), 
	.A(n2070));
   DLY4X1 FE_PHC3663_n2284 (.Y(FE_PHN3663_n2284), 
	.A(n2284));
   DLY4X1 FE_PHC3662_n2158 (.Y(FE_PHN3662_n2158), 
	.A(n2158));
   DLY4X1 FE_PHC3661_n1653 (.Y(FE_PHN3661_n1653), 
	.A(n1653));
   DLY4X1 FE_PHC3660_n1503 (.Y(FE_PHN3660_n1503), 
	.A(n1503));
   DLY4X1 FE_PHC3659_n1693 (.Y(FE_PHN3659_n1693), 
	.A(n1693));
   DLY4X1 FE_PHC3658_n2056 (.Y(FE_PHN3658_n2056), 
	.A(n2056));
   DLY4X1 FE_PHC3657_n2076 (.Y(FE_PHN3657_n2076), 
	.A(n2076));
   DLY4X1 FE_PHC3656_n1833 (.Y(FE_PHN3656_n1833), 
	.A(n1833));
   DLY4X1 FE_PHC3655_n2247 (.Y(FE_PHN3655_n2247), 
	.A(n2247));
   DLY4X1 FE_PHC3654_n1834 (.Y(FE_PHN3654_n1834), 
	.A(n1834));
   DLY4X1 FE_PHC3653_n2042 (.Y(FE_PHN3653_n2042), 
	.A(n2042));
   DLY4X1 FE_PHC3652_n1679 (.Y(FE_PHN3652_n1679), 
	.A(n1679));
   DLY4X1 FE_PHC3651_n1425 (.Y(FE_PHN3651_n1425), 
	.A(n1425));
   DLY4X1 FE_PHC3650_n1412 (.Y(FE_PHN3650_n1412), 
	.A(n1412));
   DLY4X1 FE_PHC3649_n1682 (.Y(FE_PHN3649_n1682), 
	.A(n1682));
   DLY4X1 FE_PHC3648_n1678 (.Y(FE_PHN3648_n1678), 
	.A(n1678));
   DLY4X1 FE_PHC3647_n1423 (.Y(FE_PHN3647_n1423), 
	.A(n1423));
   DLY4X1 FE_PHC3646_n1994 (.Y(FE_PHN3646_n1994), 
	.A(n1994));
   DLY4X1 FE_PHC3645_n1666 (.Y(FE_PHN3645_n1666), 
	.A(n1666));
   DLY4X1 FE_PHC3644_n2152 (.Y(FE_PHN3644_n2152), 
	.A(n2152));
   DLY4X1 FE_PHC3643_n1713 (.Y(FE_PHN3643_n1713), 
	.A(n1713));
   DLY4X1 FE_PHC3642_n2105 (.Y(FE_PHN3642_n2105), 
	.A(n2105));
   DLY4X1 FE_PHC3641_n1712 (.Y(FE_PHN3641_n1712), 
	.A(n1712));
   DLY4X1 FE_PHC3640_n2073 (.Y(FE_PHN3640_n2073), 
	.A(n2073));
   DLY4X1 FE_PHC3639_n2124 (.Y(FE_PHN3639_n2124), 
	.A(n2124));
   DLY4X1 FE_PHC3638_n1405 (.Y(FE_PHN3638_n1405), 
	.A(n1405));
   DLY4X1 FE_PHC3637_n2154 (.Y(FE_PHN3637_n2154), 
	.A(n2154));
   DLY4X1 FE_PHC3636_n2220 (.Y(FE_PHN3636_n2220), 
	.A(n2220));
   DLY4X1 FE_PHC3635_n2126 (.Y(FE_PHN3635_n2126), 
	.A(n2126));
   DLY4X1 FE_PHC3634_n1848 (.Y(FE_PHN3634_n1848), 
	.A(n1848));
   DLY4X1 FE_PHC3633_n1416 (.Y(FE_PHN3633_n1416), 
	.A(n1416));
   DLY4X1 FE_PHC3632_n2231 (.Y(FE_PHN3632_n2231), 
	.A(n2231));
   DLY4X1 FE_PHC3631_n1771 (.Y(FE_PHN3631_n1771), 
	.A(n1771));
   DLY4X1 FE_PHC3630_n1720 (.Y(FE_PHN3630_n1720), 
	.A(n1720));
   DLY4X1 FE_PHC3629_n2212 (.Y(FE_PHN3629_n2212), 
	.A(n2212));
   DLY4X1 FE_PHC3628_n2193 (.Y(FE_PHN3628_n2193), 
	.A(n2193));
   DLY4X1 FE_PHC3627_n2255 (.Y(FE_PHN3627_n2255), 
	.A(n2255));
   DLY4X1 FE_PHC3626_n2235 (.Y(FE_PHN3626_n2235), 
	.A(n2235));
   DLY4X1 FE_PHC3625_n1482 (.Y(FE_PHN3625_n1482), 
	.A(n1482));
   DLY4X1 FE_PHC3624_n2266 (.Y(FE_PHN3624_n2266), 
	.A(n2266));
   DLY4X1 FE_PHC3623_n1718 (.Y(FE_PHN3623_n1718), 
	.A(n1718));
   DLY4X1 FE_PHC3622_n1450 (.Y(FE_PHN3622_n1450), 
	.A(n1450));
   DLY4X1 FE_PHC3621_n2121 (.Y(FE_PHN3621_n2121), 
	.A(n2121));
   DLY4X1 FE_PHC3620_n1658 (.Y(FE_PHN3620_n1658), 
	.A(n1658));
   DLY4X1 FE_PHC3619_n1724 (.Y(FE_PHN3619_n1724), 
	.A(n1724));
   DLY4X1 FE_PHC3618_n2215 (.Y(FE_PHN3618_n2215), 
	.A(n2215));
   DLY4X1 FE_PHC3617_n2137 (.Y(FE_PHN3617_n2137), 
	.A(n2137));
   DLY4X1 FE_PHC3616_n1717 (.Y(FE_PHN3616_n1717), 
	.A(n1717));
   DLY4X1 FE_PHC3615_n1878 (.Y(FE_PHN3615_n1878), 
	.A(n1878));
   DLY4X1 FE_PHC3614_n1891 (.Y(FE_PHN3614_n1891), 
	.A(n1891));
   DLY4X1 FE_PHC3613_n1796 (.Y(FE_PHN3613_n1796), 
	.A(n1796));
   DLY4X1 FE_PHC3612_n1763 (.Y(FE_PHN3612_n1763), 
	.A(n1763));
   DLY4X1 FE_PHC3611_n1661 (.Y(FE_PHN3611_n1661), 
	.A(n1661));
   DLY3X1 FE_PHC3444_key_mem_1407_ (.Y(FE_PHN3444_key_mem_1407_), 
	.A(key_mem[1407]));
   DLY4X1 FE_PHC3437_key_mem_514_ (.Y(FE_PHN3437_key_mem_514_), 
	.A(key_mem[514]));
   DLY4X1 FE_PHC3435_key_mem_1299_ (.Y(FE_PHN3435_key_mem_1299_), 
	.A(key_mem[1299]));
   DLY4X1 FE_PHC3434_key_mem_898_ (.Y(FE_PHN3434_key_mem_898_), 
	.A(key_mem[898]));
   DLY4X1 FE_PHC3433_key_mem_969_ (.Y(FE_PHN3433_key_mem_969_), 
	.A(key_mem[969]));
   DLY4X1 FE_PHC3431_key_mem_1007_ (.Y(FE_PHN3431_key_mem_1007_), 
	.A(key_mem[1007]));
   DLY4X1 FE_PHC3430_key_mem_394_ (.Y(FE_PHN3430_key_mem_394_), 
	.A(key_mem[394]));
   DLY4X1 FE_PHC3429_key_mem_130_ (.Y(FE_PHN3429_key_mem_130_), 
	.A(key_mem[130]));
   DLY3X1 FE_PHC3428_key_mem_138_ (.Y(FE_PHN3428_key_mem_138_), 
	.A(key_mem[138]));
   DLY4X1 FE_PHC3427_key_mem_239_ (.Y(FE_PHN3427_key_mem_239_), 
	.A(key_mem[239]));
   DLY4X1 FE_PHC3426_key_mem_1002_ (.Y(FE_PHN3426_key_mem_1002_), 
	.A(key_mem[1002]));
   DLY4X1 FE_PHC3425_key_mem_409_ (.Y(FE_PHN3425_key_mem_409_), 
	.A(key_mem[409]));
   DLY4X1 FE_PHC3424_key_mem_201_ (.Y(FE_PHN3424_key_mem_201_), 
	.A(key_mem[201]));
   DLY4X1 FE_PHC3423_key_mem_234_ (.Y(FE_PHN3423_key_mem_234_), 
	.A(key_mem[234]));
   DLY4X1 FE_PHC3422_key_mem_490_ (.Y(FE_PHN3422_key_mem_490_), 
	.A(key_mem[490]));
   DLY4X1 FE_PHC3421_key_mem_874_ (.Y(FE_PHN3421_key_mem_874_), 
	.A(key_mem[874]));
   DLY4X1 FE_PHC3420_key_mem_143_ (.Y(FE_PHN3420_key_mem_143_), 
	.A(key_mem[143]));
   DLY4X1 FE_PHC3419_key_mem_1391_ (.Y(FE_PHN3419_key_mem_1391_), 
	.A(key_mem[1391]));
   DLY4X1 FE_PHC3418_key_mem_255_ (.Y(FE_PHN3418_key_mem_255_), 
	.A(key_mem[255]));
   DLY4X1 FE_PHC3417_key_mem_777_ (.Y(FE_PHN3417_key_mem_777_), 
	.A(key_mem[777]));
   DLY4X1 FE_PHC3416_key_mem_522_ (.Y(FE_PHN3416_key_mem_522_), 
	.A(key_mem[522]));
   DLY4X1 FE_PHC3415_key_mem_618_ (.Y(FE_PHN3415_key_mem_618_), 
	.A(key_mem[618]));
   DLY4X1 FE_PHC3414_key_mem_585_ (.Y(FE_PHN3414_key_mem_585_), 
	.A(key_mem[585]));
   DLY4X1 FE_PHC3413_key_mem_623_ (.Y(FE_PHN3413_key_mem_623_), 
	.A(key_mem[623]));
   DLY4X1 FE_PHC3412_key_mem_770_ (.Y(FE_PHN3412_key_mem_770_), 
	.A(key_mem[770]));
   DLY4X1 FE_PHC3411_key_mem_159_ (.Y(FE_PHN3411_key_mem_159_), 
	.A(key_mem[159]));
   DLY4X1 FE_PHC3410_key_mem_543_ (.Y(FE_PHN3410_key_mem_543_), 
	.A(key_mem[543]));
   CLKBUFX1 FE_PHC3409_n2430 (.Y(FE_PHN3409_n2430), 
	.A(n2430));
   DLY4X1 FE_PHC3407_n883 (.Y(FE_PHN3407_n883), 
	.A(n883));
   DLY4X1 FE_PHC3406_n881 (.Y(FE_PHN3406_n881), 
	.A(n881));
   DLY4X1 FE_PHC3403_n2427 (.Y(FE_PHN3403_n2427), 
	.A(n2427));
   DLY3X1 FE_PHC3373_n2868 (.Y(FE_PHN3373_n2868), 
	.A(n2868));
   DLY4X1 FE_PHC3319_key_mem_1183_ (.Y(FE_PHN3319_key_mem_1183_), 
	.A(key_mem[1183]));
   DLY4X1 FE_PHC3307_key_mem_1130_ (.Y(FE_PHN3307_key_mem_1130_), 
	.A(key_mem[1130]));
   DLY3X1 FE_PHC3303_key_mem_1034_ (.Y(FE_PHN3303_key_mem_1034_), 
	.A(key_mem[1034]));
   DLY4X1 FE_PHC3285_key_mem_1290_ (.Y(FE_PHN3285_key_mem_1290_), 
	.A(key_mem[1290]));
   DLY4X1 FE_PHC3283_key_mem_15_ (.Y(FE_PHN3283_key_mem_15_), 
	.A(key_mem[15]));
   DLY4X1 FE_PHC3275_key_mem_895_ (.Y(FE_PHN3275_key_mem_895_), 
	.A(key_mem[895]));
   DLY3X1 FE_PHC3270_key_mem_889_ (.Y(FE_PHN3270_key_mem_889_), 
	.A(key_mem[889]));
   DLY4X1 FE_PHC3258_key_mem_1393_ (.Y(FE_PHN3258_key_mem_1393_), 
	.A(key_mem[1393]));
   DLY4X1 FE_PHC3248_key_mem_2_ (.Y(FE_PHN3248_key_mem_2_), 
	.A(key_mem[2]));
   DLY4X1 FE_PHC3239_key_mem_1026_ (.Y(FE_PHN3239_key_mem_1026_), 
	.A(key_mem[1026]));
   DLY4X1 FE_PHC3236_key_mem_879_ (.Y(FE_PHN3236_key_mem_879_), 
	.A(key_mem[879]));
   DLY4X1 FE_PHC3234_key_mem_783_ (.Y(FE_PHN3234_key_mem_783_), 
	.A(key_mem[783]));
   DLY4X1 FE_PHC3229_key_mem_1400_ (.Y(FE_PHN3229_key_mem_1400_), 
	.A(key_mem[1400]));
   DLY4X1 FE_PHC3226_key_mem_386_ (.Y(FE_PHN3226_key_mem_386_), 
	.A(key_mem[386]));
   DLY4X1 FE_PHC3221_key_mem_511_ (.Y(FE_PHN3221_key_mem_511_), 
	.A(key_mem[511]));
   DLY4X1 FE_PHC3218_key_mem_403_ (.Y(FE_PHN3218_key_mem_403_), 
	.A(key_mem[403]));
   DLY4X1 FE_PHC3215_key_mem_746_ (.Y(FE_PHN3215_key_mem_746_), 
	.A(key_mem[746]));
   DLY4X1 FE_PHC3214_key_mem_665_ (.Y(FE_PHN3214_key_mem_665_), 
	.A(key_mem[665]));
   DLY4X1 FE_PHC3213_key_mem_495_ (.Y(FE_PHN3213_key_mem_495_), 
	.A(key_mem[495]));
   DLY4X1 FE_PHC3210_key_mem_799_ (.Y(FE_PHN3210_key_mem_799_), 
	.A(key_mem[799]));
   DLY4X1 FE_PHC3209_key_mem_407_ (.Y(FE_PHN3209_key_mem_407_), 
	.A(key_mem[407]));
   DLY4X1 FE_PHC3208_key_mem_127_ (.Y(FE_PHN3208_key_mem_127_), 
	.A(key_mem[127]));
   DLY4X1 FE_PHC3207_key_mem_856_ (.Y(FE_PHN3207_key_mem_856_), 
	.A(key_mem[856]));
   DLY4X1 FE_PHC3206_key_mem_10_ (.Y(FE_PHN3206_key_mem_10_), 
	.A(key_mem[10]));
   DLY4X1 FE_PHC3205_key_mem_1289_ (.Y(FE_PHN3205_key_mem_1289_), 
	.A(key_mem[1289]));
   DLY4X1 FE_PHC3204_key_mem_399_ (.Y(FE_PHN3204_key_mem_399_), 
	.A(key_mem[399]));
   DLY4X1 FE_PHC3203_key_mem_863_ (.Y(FE_PHN3203_key_mem_863_), 
	.A(key_mem[863]));
   DLY4X1 FE_PHC3201_key_mem_95_ (.Y(FE_PHN3201_key_mem_95_), 
	.A(key_mem[95]));
   DLY3X1 FE_PHC3198_key_mem_791_ (.Y(FE_PHN3198_key_mem_791_), 
	.A(key_mem[791]));
   DLY4X1 FE_PHC3197_key_mem_457_ (.Y(FE_PHN3197_key_mem_457_), 
	.A(key_mem[457]));
   DLY4X1 FE_PHC3196_key_mem_761_ (.Y(FE_PHN3196_key_mem_761_), 
	.A(key_mem[761]));
   DLY4X1 FE_PHC3195_key_mem_402_ (.Y(FE_PHN3195_key_mem_402_), 
	.A(key_mem[402]));
   DLY4X1 FE_PHC3194_key_mem_18_ (.Y(FE_PHN3194_key_mem_18_), 
	.A(key_mem[18]));
   DLY4X1 FE_PHC3189_key_mem_73_ (.Y(FE_PHN3189_key_mem_73_), 
	.A(key_mem[73]));
   DLY4X1 FE_PHC3188_key_mem_19_ (.Y(FE_PHN3188_key_mem_19_), 
	.A(key_mem[19]));
   DLY4X1 FE_PHC3187_key_mem_111_ (.Y(FE_PHN3187_key_mem_111_), 
	.A(key_mem[111]));
   DLY4X1 FE_PHC3186_key_mem_841_ (.Y(FE_PHN3186_key_mem_841_), 
	.A(key_mem[841]));
   DLY4X1 FE_PHC3185_key_mem_106_ (.Y(FE_PHN3185_key_mem_106_), 
	.A(key_mem[106]));
   DLY4X1 FE_PHC3184_key_mem_415_ (.Y(FE_PHN3184_key_mem_415_), 
	.A(key_mem[415]));
   DLY3X1 FE_PHC3094_key_mem_1303_ (.Y(FE_PHN3094_key_mem_1303_), 
	.A(key_mem[1303]));
   DLY4X1 FE_PHC3091_key_mem_1279_ (.Y(FE_PHN3091_key_mem_1279_), 
	.A(key_mem[1279]));
   DLY4X1 FE_PHC3089_key_mem_126_ (.Y(FE_PHN3089_key_mem_126_), 
	.A(key_mem[126]));
   DLY4X1 FE_PHC3085_key_mem_31_ (.Y(FE_PHN3085_key_mem_31_), 
	.A(key_mem[31]));
   DLY3X1 FE_PHC2855_n2423 (.Y(FE_PHN2855_n2423), 
	.A(n2423));
   DLY3X1 FE_PHC2842_key_mem_1263_ (.Y(FE_PHN2842_key_mem_1263_), 
	.A(key_mem[1263]));
   DLY4X1 FE_PHC2841_key_mem_1353_ (.Y(FE_PHN2841_key_mem_1353_), 
	.A(key_mem[1353]));
   DLY4X1 FE_PHC2840_key_mem_1295_ (.Y(FE_PHN2840_key_mem_1295_), 
	.A(key_mem[1295]));
   DLY3X1 FE_PHC2839_key_mem_1171_ (.Y(FE_PHN2839_key_mem_1171_), 
	.A(key_mem[1171]));
   DLY4X1 FE_PHC2838_key_mem_1033_ (.Y(FE_PHN2838_key_mem_1033_), 
	.A(key_mem[1033]));
   DLY4X1 FE_PHC2837_key_mem_1297_ (.Y(FE_PHN2837_key_mem_1297_), 
	.A(key_mem[1297]));
   DLY3X1 FE_PHC2836_key_mem_1382_ (.Y(FE_PHN2836_key_mem_1382_), 
	.A(key_mem[1382]));
   DLY4X1 FE_PHC2835_key_mem_1302_ (.Y(FE_PHN2835_key_mem_1302_), 
	.A(key_mem[1302]));
   DLY4X1 FE_PHC2834_key_mem_1401_ (.Y(FE_PHN2834_key_mem_1401_), 
	.A(key_mem[1401]));
   DLY4X1 FE_PHC2833_key_mem_1375_ (.Y(FE_PHN2833_key_mem_1375_), 
	.A(key_mem[1375]));
   DLY4X1 FE_PHC2832_key_mem_650_ (.Y(FE_PHN2832_key_mem_650_), 
	.A(key_mem[650]));
   DLY4X1 FE_PHC2831_key_mem_1262_ (.Y(FE_PHN2831_key_mem_1262_), 
	.A(key_mem[1262]));
   DLY4X1 FE_PHC2830_key_mem_1368_ (.Y(FE_PHN2830_key_mem_1368_), 
	.A(key_mem[1368]));
   DLY4X1 FE_PHC2829_key_mem_1305_ (.Y(FE_PHN2829_key_mem_1305_), 
	.A(key_mem[1305]));
   DLY4X1 FE_PHC2828_key_mem_1351_ (.Y(FE_PHN2828_key_mem_1351_), 
	.A(key_mem[1351]));
   DLY4X1 FE_PHC2827_key_mem_1304_ (.Y(FE_PHN2827_key_mem_1304_), 
	.A(key_mem[1304]));
   DLY4X1 FE_PHC2826_key_mem_504_ (.Y(FE_PHN2826_key_mem_504_), 
	.A(key_mem[504]));
   DLY4X1 FE_PHC2825_key_mem_1282_ (.Y(FE_PHN2825_key_mem_1282_), 
	.A(key_mem[1282]));
   DLY4X1 FE_PHC2824_key_mem_753_ (.Y(FE_PHN2824_key_mem_753_), 
	.A(key_mem[753]));
   DLY4X1 FE_PHC2823_key_mem_1298_ (.Y(FE_PHN2823_key_mem_1298_), 
	.A(key_mem[1298]));
   DLY2X1 FE_PHC2820_n2421 (.Y(FE_PHN2820_n2421), 
	.A(n2421));
   DLY2X1 FE_PHC2814_n880 (.Y(FE_PHN2814_n880), 
	.A(n880));
   DLY3X1 FE_PHC2811_n2422 (.Y(FE_PHN2811_n2422), 
	.A(n2422));
   DLY4X1 FE_PHC2810_key_mem_1386_ (.Y(FE_PHN2810_key_mem_1386_), 
	.A(key_mem[1386]));
   DLY4X1 FE_PHC2799_n2391 (.Y(FE_PHN2799_n2391), 
	.A(FE_PHN5061_n2391));
   DLY4X1 FE_PHC2798_n2392 (.Y(FE_PHN2798_n2392), 
	.A(FE_PHN5058_n2392));
   DLY4X1 FE_PHC2795_n2390 (.Y(FE_PHN2795_n2390), 
	.A(FE_PHN5032_n2390));
   DLY4X1 FE_PHC2793_n2396 (.Y(FE_PHN2793_n2396), 
	.A(FE_PHN5027_n2396));
   DLY4X1 FE_PHC2792_n2395 (.Y(FE_PHN2792_n2395), 
	.A(FE_PHN5020_n2395));
   DLY4X1 FE_PHC2791_n2389 (.Y(FE_PHN2791_n2389), 
	.A(FE_PHN4997_n2389));
   DLY4X1 FE_PHC2790_n957 (.Y(FE_PHN2790_n957), 
	.A(FE_PHN4970_n957));
   DLY4X1 FE_PHC2789_key_mem_846_ (.Y(FE_PHN2789_key_mem_846_), 
	.A(FE_PHN4996_key_mem_846_));
   DLY4X1 FE_PHC2788_n918 (.Y(FE_PHN2788_n918), 
	.A(FE_PHN4965_n918));
   DLY4X1 FE_PHC2787_n1230 (.Y(FE_PHN2787_n1230), 
	.A(FE_PHN4855_n1230));
   DLY4X1 FE_PHC2786_n992 (.Y(FE_PHN2786_n992), 
	.A(FE_PHN4938_n992));
   DLY4X1 FE_PHC2785_n1329 (.Y(FE_PHN2785_n1329), 
	.A(FE_PHN4977_n1329));
   DLY4X1 FE_PHC2784_n935 (.Y(FE_PHN2784_n935), 
	.A(FE_PHN4859_n935));
   DLY4X1 FE_PHC2783_n1348 (.Y(FE_PHN2783_n1348), 
	.A(FE_PHN4817_n1348));
   DLY4X1 FE_PHC2782_n1355 (.Y(FE_PHN2782_n1355), 
	.A(FE_PHN4813_n1355));
   DLY4X1 FE_PHC2781_n1393 (.Y(FE_PHN2781_n1393), 
	.A(FE_PHN4867_n1393));
   DLY4X1 FE_PHC2780_n1371 (.Y(FE_PHN2780_n1371), 
	.A(FE_PHN4887_n1371));
   DLY4X1 FE_PHC2779_n965 (.Y(FE_PHN2779_n965), 
	.A(FE_PHN4939_n965));
   DLY4X1 FE_PHC2778_n973 (.Y(FE_PHN2778_n973), 
	.A(FE_PHN4732_n973));
   DLY4X1 FE_PHC2777_n886 (.Y(FE_PHN2777_n886), 
	.A(FE_PHN4871_n886));
   DLY4X1 FE_PHC2776_n1344 (.Y(FE_PHN2776_n1344), 
	.A(FE_PHN4872_n1344));
   DLY4X1 FE_PHC2775_n1294 (.Y(FE_PHN2775_n1294), 
	.A(FE_PHN4780_n1294));
   DLY4X1 FE_PHC2774_n1357 (.Y(FE_PHN2774_n1357), 
	.A(FE_PHN4793_n1357));
   DLY4X1 FE_PHC2773_n1319 (.Y(FE_PHN2773_n1319), 
	.A(FE_PHN4956_n1319));
   DLY4X1 FE_PHC2772_n931 (.Y(FE_PHN2772_n931), 
	.A(FE_PHN4952_n931));
   DLY4X1 FE_PHC2771_n1390 (.Y(FE_PHN2771_n1390), 
	.A(FE_PHN4955_n1390));
   DLY4X1 FE_PHC2770_n974 (.Y(FE_PHN2770_n974), 
	.A(FE_PHN4897_n974));
   DLY4X1 FE_PHC2769_n1075 (.Y(FE_PHN2769_n1075), 
	.A(FE_PHN4719_n1075));
   DLY4X1 FE_PHC2768_n1338 (.Y(FE_PHN2768_n1338), 
	.A(FE_PHN4727_n1338));
   DLY4X1 FE_PHC2767_n958 (.Y(FE_PHN2767_n958), 
	.A(FE_PHN4896_n958));
   DLY4X1 FE_PHC2766_n1363 (.Y(FE_PHN2766_n1363), 
	.A(FE_PHN4641_n1363));
   DLY4X1 FE_PHC2765_n1332 (.Y(FE_PHN2765_n1332), 
	.A(FE_PHN4590_n1332));
   DLY4X1 FE_PHC2764_n1380 (.Y(FE_PHN2764_n1380), 
	.A(FE_PHN4599_n1380));
   DLY4X1 FE_PHC2763_n1361 (.Y(FE_PHN2763_n1361), 
	.A(FE_PHN4549_n1361));
   DLY4X1 FE_PHC2762_n1356 (.Y(FE_PHN2762_n1356), 
	.A(FE_PHN4865_n1356));
   DLY4X1 FE_PHC2761_n1008 (.Y(FE_PHN2761_n1008), 
	.A(FE_PHN4499_n1008));
   DLY4X1 FE_PHC2760_n1387 (.Y(FE_PHN2760_n1387), 
	.A(FE_PHN4593_n1387));
   DLY4X1 FE_PHC2759_n1009 (.Y(FE_PHN2759_n1009), 
	.A(FE_PHN4847_n1009));
   DLY4X1 FE_PHC2758_n997 (.Y(FE_PHN2758_n997), 
	.A(n997));
   DLY4X1 FE_PHC2757_n954 (.Y(FE_PHN2757_n954), 
	.A(FE_PHN4827_n954));
   DLY4X1 FE_PHC2756_n2188 (.Y(FE_PHN2756_n2188), 
	.A(FE_PHN4731_n2188));
   DLY4X1 FE_PHC2755_n2091 (.Y(FE_PHN2755_n2091), 
	.A(n2091));
   DLY4X1 FE_PHC2754_n926 (.Y(FE_PHN2754_n926), 
	.A(FE_PHN4756_n926));
   DLY4X1 FE_PHC2753_n2229 (.Y(FE_PHN2753_n2229), 
	.A(FE_PHN4885_n2229));
   DLY4X1 FE_PHC2752_n1327 (.Y(FE_PHN2752_n1327), 
	.A(FE_PHN4945_n1327));
   DLY4X1 FE_PHC2751_n1340 (.Y(FE_PHN2751_n1340), 
	.A(FE_PHN4317_n1340));
   DLY4X1 FE_PHC2750_n1879 (.Y(FE_PHN2750_n1879), 
	.A(FE_PHN4517_n1879));
   DLY4X1 FE_PHC2749_n1298 (.Y(FE_PHN2749_n1298), 
	.A(FE_PHN4405_n1298));
   DLY4X1 FE_PHC2748_n1284 (.Y(FE_PHN2748_n1284), 
	.A(FE_PHN4714_n1284));
   DLY4X1 FE_PHC2747_n1744 (.Y(FE_PHN2747_n1744), 
	.A(n1744));
   DLY4X1 FE_PHC2746_n1856 (.Y(FE_PHN2746_n1856), 
	.A(FE_PHN4472_n1856));
   DLY4X1 FE_PHC2745_n1272 (.Y(FE_PHN2745_n1272), 
	.A(FE_PHN4626_n1272));
   DLY4X1 FE_PHC2744_n1359 (.Y(FE_PHN2744_n1359), 
	.A(FE_PHN4947_n1359));
   DLY4X1 FE_PHC2743_n1368 (.Y(FE_PHN2743_n1368), 
	.A(FE_PHN4398_n1368));
   DLY4X1 FE_PHC2742_n932 (.Y(FE_PHN2742_n932), 
	.A(FE_PHN4628_n932));
   DLY4X1 FE_PHC2741_n1350 (.Y(FE_PHN2741_n1350), 
	.A(FE_PHN4702_n1350));
   DLY4X1 FE_PHC2740_n942 (.Y(FE_PHN2740_n942), 
	.A(FE_PHN4466_n942));
   DLY4X1 FE_PHC2739_n1339 (.Y(FE_PHN2739_n1339), 
	.A(FE_PHN4687_n1339));
   DLY4X1 FE_PHC2738_n885 (.Y(FE_PHN2738_n885), 
	.A(n885));
   DLY4X1 FE_PHC2737_n1276 (.Y(FE_PHN2737_n1276), 
	.A(FE_PHN4761_n1276));
   DLY4X1 FE_PHC2736_n1269 (.Y(FE_PHN2736_n1269), 
	.A(FE_PHN4441_n1269));
   DLY4X1 FE_PHC2735_n1351 (.Y(FE_PHN2735_n1351), 
	.A(FE_PHN4363_n1351));
   DLY4X1 FE_PHC2734_n1286 (.Y(FE_PHN2734_n1286), 
	.A(FE_PHN4416_n1286));
   DLY4X1 FE_PHC2733_n1352 (.Y(FE_PHN2733_n1352), 
	.A(FE_PHN4643_n1352));
   DLY4X1 FE_PHC2732_n1315 (.Y(FE_PHN2732_n1315), 
	.A(FE_PHN4674_n1315));
   DLY4X1 FE_PHC2731_n939 (.Y(FE_PHN2731_n939), 
	.A(n939));
   DLY4X1 FE_PHC2730_n1005 (.Y(FE_PHN2730_n1005), 
	.A(FE_PHN4556_n1005));
   DLY4X1 FE_PHC2729_n1307 (.Y(FE_PHN2729_n1307), 
	.A(FE_PHN4801_n1307));
   DLY4X1 FE_PHC2728_n2149 (.Y(FE_PHN2728_n2149), 
	.A(FE_PHN4449_n2149));
   DLY4X1 FE_PHC2727_n1501 (.Y(FE_PHN2727_n1501), 
	.A(n1501));
   DLY4X1 FE_PHC2726_n1349 (.Y(FE_PHN2726_n1349), 
	.A(FE_PHN4743_n1349));
   DLY4X1 FE_PHC2725_n1384 (.Y(FE_PHN2725_n1384), 
	.A(FE_PHN4456_n1384));
   DLY4X1 FE_PHC2724_n1301 (.Y(FE_PHN2724_n1301), 
	.A(FE_PHN4321_n1301));
   DLY4X1 FE_PHC2723_n925 (.Y(FE_PHN2723_n925), 
	.A(FE_PHN4671_n925));
   DLY4X1 FE_PHC2722_n963 (.Y(FE_PHN2722_n963), 
	.A(FE_PHN4382_n963));
   DLY4X1 FE_PHC2721_n960 (.Y(FE_PHN2721_n960), 
	.A(FE_PHN4597_n960));
   DLY4X1 FE_PHC2720_n977 (.Y(FE_PHN2720_n977), 
	.A(FE_PHN4596_n977));
   DLY4X1 FE_PHC2719_n1358 (.Y(FE_PHN2719_n1358), 
	.A(FE_PHN4535_n1358));
   DLY4X1 FE_PHC2718_n1303 (.Y(FE_PHN2718_n1303), 
	.A(FE_PHN4678_n1303));
   DLY4X1 FE_PHC2717_n1468 (.Y(FE_PHN2717_n1468), 
	.A(FE_PHN4511_n1468));
   DLY4X1 FE_PHC2716_n1812 (.Y(FE_PHN2716_n1812), 
	.A(FE_PHN4577_n1812));
   DLY4X1 FE_PHC2715_n1392 (.Y(FE_PHN2715_n1392), 
	.A(FE_PHN4682_n1392));
   DLY4X1 FE_PHC2714_n1378 (.Y(FE_PHN2714_n1378), 
	.A(FE_PHN4423_n1378));
   DLY4X1 FE_PHC2713_n928 (.Y(FE_PHN2713_n928), 
	.A(FE_PHN4483_n928));
   DLY4X1 FE_PHC2712_n1001 (.Y(FE_PHN2712_n1001), 
	.A(FE_PHN4880_n1001));
   DLY4X1 FE_PHC2711_n1853 (.Y(FE_PHN2711_n1853), 
	.A(FE_PHN4420_n1853));
   DLY4X1 FE_PHC2710_n1278 (.Y(FE_PHN2710_n1278), 
	.A(FE_PHN4503_n1278));
   DLY4X1 FE_PHC2709_n1275 (.Y(FE_PHN2709_n1275), 
	.A(FE_PHN4341_n1275));
   DLY4X1 FE_PHC2708_n1377 (.Y(FE_PHN2708_n1377), 
	.A(FE_PHN4361_n1377));
   DLY4X1 FE_PHC2707_n2114 (.Y(FE_PHN2707_n2114), 
	.A(n2114));
   DLY4X1 FE_PHC2706_n1341 (.Y(FE_PHN2706_n1341), 
	.A(FE_PHN4510_n1341));
   DLY4X1 FE_PHC2705_n1839 (.Y(FE_PHN2705_n1839), 
	.A(FE_PHN4237_n1839));
   DLY4X1 FE_PHC2704_n1293 (.Y(FE_PHN2704_n1293), 
	.A(FE_PHN4886_n1293));
   DLY4X1 FE_PHC2703_n993 (.Y(FE_PHN2703_n993), 
	.A(n993));
   DLY4X1 FE_PHC2702_n899 (.Y(FE_PHN2702_n899), 
	.A(n899));
   DLY4X1 FE_PHC2701_n1886 (.Y(FE_PHN2701_n1886), 
	.A(FE_PHN4901_n1886));
   DLY4X1 FE_PHC2700_n887 (.Y(FE_PHN2700_n887), 
	.A(FE_PHN4612_n887));
   DLY4X1 FE_PHC2699_n1372 (.Y(FE_PHN2699_n1372), 
	.A(FE_PHN4324_n1372));
   DLY4X1 FE_PHC2698_n937 (.Y(FE_PHN2698_n937), 
	.A(FE_PHN4125_n937));
   DLY4X1 FE_PHC2697_n2180 (.Y(FE_PHN2697_n2180), 
	.A(FE_PHN4730_n2180));
   DLY4X1 FE_PHC2696_n1109 (.Y(FE_PHN2696_n1109), 
	.A(n1109));
   DLY4X1 FE_PHC2695_n1790 (.Y(FE_PHN2695_n1790), 
	.A(FE_PHN4293_n1790));
   DLY4X1 FE_PHC2694_n1292 (.Y(FE_PHN2694_n1292), 
	.A(FE_PHN4390_n1292));
   DLY4X1 FE_PHC2693_n2046 (.Y(FE_PHN2693_n2046), 
	.A(n2046));
   DLY4X1 FE_PHC2692_n995 (.Y(FE_PHN2692_n995), 
	.A(n995));
   DLY4X1 FE_PHC2691_n1302 (.Y(FE_PHN2691_n1302), 
	.A(FE_PHN4763_n1302));
   DLY4X1 FE_PHC2690_n915 (.Y(FE_PHN2690_n915), 
	.A(FE_PHN4709_n915));
   DLY4X1 FE_PHC2689_n1867 (.Y(FE_PHN2689_n1867), 
	.A(n1867));
   DLY4X1 FE_PHC2688_n1330 (.Y(FE_PHN2688_n1330), 
	.A(FE_PHN4150_n1330));
   DLY4X1 FE_PHC2687_n1007 (.Y(FE_PHN2687_n1007), 
	.A(FE_PHN4618_n1007));
   DLY4X1 FE_PHC2686_n1383 (.Y(FE_PHN2686_n1383), 
	.A(FE_PHN4560_n1383));
   DLY4X1 FE_PHC2685_n999 (.Y(FE_PHN2685_n999), 
	.A(FE_PHN4554_n999));
   DLY4X1 FE_PHC2684_n929 (.Y(FE_PHN2684_n929), 
	.A(FE_PHN4325_n929));
   DLY4X1 FE_PHC2683_n1375 (.Y(FE_PHN2683_n1375), 
	.A(FE_PHN4181_n1375));
   DLY4X1 FE_PHC2682_n1432 (.Y(FE_PHN2682_n1432), 
	.A(FE_PHN4428_n1432));
   DLY4X1 FE_PHC2681_n1311 (.Y(FE_PHN2681_n1311), 
	.A(FE_PHN4185_n1311));
   DLY4X1 FE_PHC2680_n1346 (.Y(FE_PHN2680_n1346), 
	.A(FE_PHN4309_n1346));
   DLY4X1 FE_PHC2679_n1872 (.Y(FE_PHN2679_n1872), 
	.A(FE_PHN4839_n1872));
   DLY4X1 FE_PHC2678_n1281 (.Y(FE_PHN2678_n1281), 
	.A(FE_PHN4615_n1281));
   DLY4X1 FE_PHC2677_n2116 (.Y(FE_PHN2677_n2116), 
	.A(FE_PHN4657_n2116));
   DLY4X1 FE_PHC2676_n1836 (.Y(FE_PHN2676_n1836), 
	.A(FE_PHN4623_n1836));
   DLY4X1 FE_PHC2675_n896 (.Y(FE_PHN2675_n896), 
	.A(FE_PHN4467_n896));
   DLY4X1 FE_PHC2674_n1002 (.Y(FE_PHN2674_n1002), 
	.A(n1002));
   DLY4X1 FE_PHC2673_n1347 (.Y(FE_PHN2673_n1347), 
	.A(FE_PHN4241_n1347));
   DLY4X1 FE_PHC2672_n1374 (.Y(FE_PHN2672_n1374), 
	.A(FE_PHN4415_n1374));
   DLY4X1 FE_PHC2671_n1493 (.Y(FE_PHN2671_n1493), 
	.A(n1493));
   DLY4X1 FE_PHC2670_n2228 (.Y(FE_PHN2670_n2228), 
	.A(n2228));
   DLY4X1 FE_PHC2669_n1765 (.Y(FE_PHN2669_n1765), 
	.A(FE_PHN4228_n1765));
   DLY4X1 FE_PHC2668_n2045 (.Y(FE_PHN2668_n2045), 
	.A(FE_PHN4236_n2045));
   DLY4X1 FE_PHC2667_n2119 (.Y(FE_PHN2667_n2119), 
	.A(FE_PHN4634_n2119));
   DLY4X1 FE_PHC2666_n1337 (.Y(FE_PHN2666_n1337), 
	.A(FE_PHN4103_n1337));
   DLY4X1 FE_PHC2665_n986 (.Y(FE_PHN2665_n986), 
	.A(FE_PHN4024_n986));
   DLY4X1 FE_PHC2664_n1746 (.Y(FE_PHN2664_n1746), 
	.A(FE_PHN4684_n1746));
   DLY4X1 FE_PHC2663_n1270 (.Y(FE_PHN2663_n1270), 
	.A(FE_PHN4454_n1270));
   DLY4X1 FE_PHC2662_n919 (.Y(FE_PHN2662_n919), 
	.A(FE_PHN4213_n919));
   DLY4X1 FE_PHC2661_n1810 (.Y(FE_PHN2661_n1810), 
	.A(FE_PHN4360_n1810));
   DLY4X1 FE_PHC2660_n998 (.Y(FE_PHN2660_n998), 
	.A(FE_PHN4370_n998));
   DLY4X1 FE_PHC2659_n1430 (.Y(FE_PHN2659_n1430), 
	.A(FE_PHN4175_n1430));
   DLY4X1 FE_PHC2658_n2060 (.Y(FE_PHN2658_n2060), 
	.A(FE_PHN4676_n2060));
   DLY4X1 FE_PHC2657_n914 (.Y(FE_PHN2657_n914), 
	.A(FE_PHN4494_n914));
   DLY4X1 FE_PHC2656_n1322 (.Y(FE_PHN2656_n1322), 
	.A(FE_PHN4660_n1322));
   DLY4X1 FE_PHC2655_n2038 (.Y(FE_PHN2655_n2038), 
	.A(FE_PHN4180_n2038));
   DLY4X1 FE_PHC2654_n1408 (.Y(FE_PHN2654_n1408), 
	.A(n1408));
   DLY4X1 FE_PHC2653_n1324 (.Y(FE_PHN2653_n1324), 
	.A(FE_PHN4661_n1324));
   DLY4X1 FE_PHC2652_n940 (.Y(FE_PHN2652_n940), 
	.A(FE_PHN4127_n940));
   DLY4X1 FE_PHC2651_n1388 (.Y(FE_PHN2651_n1388), 
	.A(FE_PHN4595_n1388));
   DLY4X1 FE_PHC2650_n1479 (.Y(FE_PHN2650_n1479), 
	.A(FE_PHN4344_n1479));
   DLY4X1 FE_PHC2649_n2111 (.Y(FE_PHN2649_n2111), 
	.A(FE_PHN4273_n2111));
   DLY4X1 FE_PHC2648_n1516 (.Y(FE_PHN2648_n1516), 
	.A(FE_PHN4214_n1516));
   DLY4X1 FE_PHC2647_n1312 (.Y(FE_PHN2647_n1312), 
	.A(FE_PHN4473_n1312));
   DLY4X1 FE_PHC2646_n1271 (.Y(FE_PHN2646_n1271), 
	.A(FE_PHN4080_n1271));
   DLY4X1 FE_PHC2645_n2189 (.Y(FE_PHN2645_n2189), 
	.A(n2189));
   DLY4X1 FE_PHC2644_n1427 (.Y(FE_PHN2644_n1427), 
	.A(FE_PHN4159_n1427));
   DLY4X1 FE_PHC2643_n1304 (.Y(FE_PHN2643_n1304), 
	.A(FE_PHN4857_n1304));
   DLY4X1 FE_PHC2642_n1784 (.Y(FE_PHN2642_n1784), 
	.A(FE_PHN4238_n1784));
   DLY4X1 FE_PHC2641_n907 (.Y(FE_PHN2641_n907), 
	.A(FE_PHN4614_n907));
   DLY4X1 FE_PHC2640_n989 (.Y(FE_PHN2640_n989), 
	.A(n989));
   DLY4X1 FE_PHC2639_n1289 (.Y(FE_PHN2639_n1289), 
	.A(FE_PHN4373_n1289));
   DLY4X1 FE_PHC2638_n1758 (.Y(FE_PHN2638_n1758), 
	.A(n1758));
   DLY4X1 FE_PHC2637_n1775 (.Y(FE_PHN2637_n1775), 
	.A(FE_PHN4114_n1775));
   DLY4X1 FE_PHC2636_n2234 (.Y(FE_PHN2636_n2234), 
	.A(FE_PHN4408_n2234));
   DLY4X1 FE_PHC2635_n1749 (.Y(FE_PHN2635_n1749), 
	.A(FE_PHN4386_n1749));
   DLY4X1 FE_PHC2634_n894 (.Y(FE_PHN2634_n894), 
	.A(FE_PHN4003_n894));
   DLY4X1 FE_PHC2633_n956 (.Y(FE_PHN2633_n956), 
	.A(FE_PHN4409_n956));
   DLY4X1 FE_PHC2632_n1277 (.Y(FE_PHN2632_n1277), 
	.A(FE_PHN4276_n1277));
   DLY4X1 FE_PHC2631_n1333 (.Y(FE_PHN2631_n1333), 
	.A(FE_PHN4087_n1333));
   DLY4X1 FE_PHC2630_n903 (.Y(FE_PHN2630_n903), 
	.A(FE_PHN3977_n903));
   DLY4X1 FE_PHC2629_n927 (.Y(FE_PHN2629_n927), 
	.A(FE_PHN4481_n927));
   DLY4X1 FE_PHC2628_n2249 (.Y(FE_PHN2628_n2249), 
	.A(FE_PHN3931_n2249));
   DLY4X1 FE_PHC2627_n1464 (.Y(FE_PHN2627_n1464), 
	.A(FE_PHN4380_n1464));
   DLY4X1 FE_PHC2626_n2223 (.Y(FE_PHN2626_n2223), 
	.A(FE_PHN4665_n2223));
   DLY4X1 FE_PHC2625_n1522 (.Y(FE_PHN2625_n1522), 
	.A(FE_PHN4006_n1522));
   DLY4X1 FE_PHC2624_n1300 (.Y(FE_PHN2624_n1300), 
	.A(FE_PHN4805_n1300));
   DLY4X1 FE_PHC2623_n1370 (.Y(FE_PHN2623_n1370), 
	.A(FE_PHN4247_n1370));
   DLY4X1 FE_PHC2622_n1813 (.Y(FE_PHN2622_n1813), 
	.A(FE_PHN4427_n1813));
   DLY4X1 FE_PHC2621_n2290 (.Y(FE_PHN2621_n2290), 
	.A(n2290));
   DLY4X1 FE_PHC2620_n1888 (.Y(FE_PHN2620_n1888), 
	.A(FE_PHN4910_n1888));
   DLY4X1 FE_PHC2619_n1325 (.Y(FE_PHN2619_n1325), 
	.A(FE_PHN4482_n1325));
   DLY4X1 FE_PHC2618_n1517 (.Y(FE_PHN2618_n1517), 
	.A(n1517));
   DLY4X1 FE_PHC2617_n1843 (.Y(FE_PHN2617_n1843), 
	.A(n1843));
   DLY4X1 FE_PHC2616_n916 (.Y(FE_PHN2616_n916), 
	.A(FE_PHN4277_n916));
   DLY4X1 FE_PHC2615_n1309 (.Y(FE_PHN2615_n1309), 
	.A(FE_PHN4165_n1309));
   DLY4X1 FE_PHC2614_n945 (.Y(FE_PHN2614_n945), 
	.A(FE_PHN4430_n945));
   DLY4X1 FE_PHC2613_n1382 (.Y(FE_PHN2613_n1382), 
	.A(FE_PHN4002_n1382));
   DLY4X1 FE_PHC2612_n1663 (.Y(FE_PHN2612_n1663), 
	.A(FE_PHN4314_n1663));
   DLY4X1 FE_PHC2611_n1445 (.Y(FE_PHN2611_n1445), 
	.A(FE_PHN4244_n1445));
   DLY4X1 FE_PHC2610_n1291 (.Y(FE_PHN2610_n1291), 
	.A(FE_PHN4281_n1291));
   DLY4X1 FE_PHC2609_n911 (.Y(FE_PHN2609_n911), 
	.A(FE_PHN4212_n911));
   DLY4X1 FE_PHC2608_n2182 (.Y(FE_PHN2608_n2182), 
	.A(FE_PHN4547_n2182));
   DLY4X1 FE_PHC2607_n1859 (.Y(FE_PHN2607_n1859), 
	.A(FE_PHN4323_n1859));
   DLY4X1 FE_PHC2606_n1403 (.Y(FE_PHN2606_n1403), 
	.A(FE_PHN4031_n1403));
   DLY4X1 FE_PHC2605_n959 (.Y(FE_PHN2605_n959), 
	.A(FE_PHN4229_n959));
   DLY4X1 FE_PHC2604_n2287 (.Y(FE_PHN2604_n2287), 
	.A(n2287));
   DLY4X1 FE_PHC2603_n1477 (.Y(FE_PHN2603_n1477), 
	.A(FE_PHN4300_n1477));
   DLY4X1 FE_PHC2602_n983 (.Y(FE_PHN2602_n983), 
	.A(FE_PHN4395_n983));
   DLY4X1 FE_PHC2601_n1816 (.Y(FE_PHN2601_n1816), 
	.A(FE_PHN4282_n1816));
   DLY4X1 FE_PHC2600_n2065 (.Y(FE_PHN2600_n2065), 
	.A(FE_PHN4284_n2065));
   DLY4X1 FE_PHC2599_n961 (.Y(FE_PHN2599_n961), 
	.A(FE_PHN4319_n961));
   DLY4X1 FE_PHC2598_n2039 (.Y(FE_PHN2598_n2039), 
	.A(FE_PHN4095_n2039));
   DLY4X1 FE_PHC2597_n2241 (.Y(FE_PHN2597_n2241), 
	.A(FE_PHN4156_n2241));
   DLY4X1 FE_PHC2596_n1793 (.Y(FE_PHN2596_n1793), 
	.A(n1793));
   DLY4X1 FE_PHC2595_n1313 (.Y(FE_PHN2595_n1313), 
	.A(FE_PHN4620_n1313));
   DLY4X1 FE_PHC2594_n1316 (.Y(FE_PHN2594_n1316), 
	.A(FE_PHN3947_n1316));
   DLY4X1 FE_PHC2593_n1321 (.Y(FE_PHN2593_n1321), 
	.A(FE_PHN4636_n1321));
   DLY4X1 FE_PHC2592_n1455 (.Y(FE_PHN2592_n1455), 
	.A(FE_PHN4174_n1455));
   DLY4X1 FE_PHC2591_n1518 (.Y(FE_PHN2591_n1518), 
	.A(FE_PHN4122_n1518));
   DLY4X1 FE_PHC2590_n936 (.Y(FE_PHN2590_n936), 
	.A(FE_PHN4662_n936));
   DLY4X1 FE_PHC2589_n930 (.Y(FE_PHN2589_n930), 
	.A(FE_PHN3927_n930));
   DLY4X1 FE_PHC2588_n1394 (.Y(FE_PHN2588_n1394), 
	.A(n1394));
   DLY4X1 FE_PHC2587_n910 (.Y(FE_PHN2587_n910), 
	.A(n910));
   DLY4X1 FE_PHC2586_n1273 (.Y(FE_PHN2586_n1273), 
	.A(FE_PHN4096_n1273));
   DLY4X1 FE_PHC2585_n2109 (.Y(FE_PHN2585_n2109), 
	.A(FE_PHN3935_n2109));
   DLY4X1 FE_PHC2584_n1285 (.Y(FE_PHN2584_n1285), 
	.A(n1285));
   DLY4X1 FE_PHC2583_n1279 (.Y(FE_PHN2583_n1279), 
	.A(FE_PHN4275_n1279));
   DLY4X1 FE_PHC2582_n1730 (.Y(FE_PHN2582_n1730), 
	.A(FE_PHN4988_n1730));
   DLY4X1 FE_PHC2581_n900 (.Y(FE_PHN2581_n900), 
	.A(FE_PHN4303_n900));
   DLY4X1 FE_PHC2580_n1369 (.Y(FE_PHN2580_n1369), 
	.A(FE_PHN3850_n1369));
   DLY4X1 FE_PHC2579_n2271 (.Y(FE_PHN2579_n2271), 
	.A(FE_PHN4274_n2271));
   DLY4X1 FE_PHC2578_n1435 (.Y(FE_PHN2578_n1435), 
	.A(FE_PHN4094_n1435));
   DLY4X1 FE_PHC2577_n1428 (.Y(FE_PHN2577_n1428), 
	.A(FE_PHN3911_n1428));
   DLY4X1 FE_PHC2576_n2176 (.Y(FE_PHN2576_n2176), 
	.A(FE_PHN4067_n2176));
   DLY4X1 FE_PHC2575_n1716 (.Y(FE_PHN2575_n1716), 
	.A(FE_PHN4119_n1716));
   DLY4X1 FE_PHC2574_n1362 (.Y(FE_PHN2574_n1362), 
	.A(FE_PHN4308_n1362));
   DLY4X1 FE_PHC2573_n2289 (.Y(FE_PHN2573_n2289), 
	.A(FE_PHN4135_n2289));
   DLY4X1 FE_PHC2572_n1676 (.Y(FE_PHN2572_n1676), 
	.A(FE_PHN4173_n1676));
   DLY4X1 FE_PHC2571_n1449 (.Y(FE_PHN2571_n1449), 
	.A(FE_PHN4142_n1449));
   DLY4X1 FE_PHC2570_n984 (.Y(FE_PHN2570_n984), 
	.A(FE_PHN4134_n984));
   DLY4X1 FE_PHC2569_n1700 (.Y(FE_PHN2569_n1700), 
	.A(FE_PHN4288_n1700));
   DLY4X1 FE_PHC2568_n949 (.Y(FE_PHN2568_n949), 
	.A(FE_PHN4001_n949));
   DLY4X1 FE_PHC2567_n1287 (.Y(FE_PHN2567_n1287), 
	.A(FE_PHN4371_n1287));
   DLY4X1 FE_PHC2566_n2166 (.Y(FE_PHN2566_n2166), 
	.A(n2166));
   DLY4X1 FE_PHC2565_n943 (.Y(FE_PHN2565_n943), 
	.A(FE_PHN4525_n943));
   DLY4X1 FE_PHC2564_n970 (.Y(FE_PHN2564_n970), 
	.A(FE_PHN4192_n970));
   DLY4X1 FE_PHC2563_n934 (.Y(FE_PHN2563_n934), 
	.A(FE_PHN4256_n934));
   DLY4X1 FE_PHC2562_n1515 (.Y(FE_PHN2562_n1515), 
	.A(FE_PHN4038_n1515));
   DLY4X1 FE_PHC2561_n2094 (.Y(FE_PHN2561_n2094), 
	.A(FE_PHN4537_n2094));
   DLY4X1 FE_PHC2560_n2117 (.Y(FE_PHN2560_n2117), 
	.A(FE_PHN4705_n2117));
   DLY4X1 FE_PHC2559_n1689 (.Y(FE_PHN2559_n1689), 
	.A(FE_PHN4698_n1689));
   DLY4X1 FE_PHC2558_n1471 (.Y(FE_PHN2558_n1471), 
	.A(FE_PHN4085_n1471));
   DLY4X1 FE_PHC2557_n1353 (.Y(FE_PHN2557_n1353), 
	.A(FE_PHN4108_n1353));
   DLY4X1 FE_PHC2556_n988 (.Y(FE_PHN2556_n988), 
	.A(n988));
   DLY4X1 FE_PHC2555_n933 (.Y(FE_PHN2555_n933), 
	.A(FE_PHN4146_n933));
   DLY4X1 FE_PHC2554_n1400 (.Y(FE_PHN2554_n1400), 
	.A(FE_PHN3975_n1400));
   DLY4X1 FE_PHC2553_n2084 (.Y(FE_PHN2553_n2084), 
	.A(FE_PHN4734_n2084));
   DLY4X1 FE_PHC2552_n2291 (.Y(FE_PHN2552_n2291), 
	.A(FE_PHN4091_n2291));
   DLY4X1 FE_PHC2551_n909 (.Y(FE_PHN2551_n909), 
	.A(FE_PHN4607_n909));
   DLY4X1 FE_PHC2550_n1838 (.Y(FE_PHN2550_n1838), 
	.A(FE_PHN4406_n1838));
   DLY4X1 FE_PHC2549_n1402 (.Y(FE_PHN2549_n1402), 
	.A(FE_PHN3973_n1402));
   DLY4X1 FE_PHC2548_n1011 (.Y(FE_PHN2548_n1011), 
	.A(FE_PHN4149_n1011));
   DLY4X1 FE_PHC2547_n2066 (.Y(FE_PHN2547_n2066), 
	.A(FE_PHN3991_n2066));
   DLY4X1 FE_PHC2546_n1703 (.Y(FE_PHN2546_n1703), 
	.A(FE_PHN3902_n1703));
   DLY4X1 FE_PHC2545_n905 (.Y(FE_PHN2545_n905), 
	.A(FE_PHN3963_n905));
   DLY4X1 FE_PHC2544_n1500 (.Y(FE_PHN2544_n1500), 
	.A(FE_PHN4157_n1500));
   DLY4X1 FE_PHC2543_n1874 (.Y(FE_PHN2543_n1874), 
	.A(FE_PHN3894_n1874));
   DLY4X1 FE_PHC2542_n1431 (.Y(FE_PHN2542_n1431), 
	.A(FE_PHN3910_n1431));
   DLY4X1 FE_PHC2541_n1708 (.Y(FE_PHN2541_n1708), 
	.A(FE_PHN4086_n1708));
   DLY4X1 FE_PHC2540_n967 (.Y(FE_PHN2540_n967), 
	.A(FE_PHN3919_n967));
   DLY4X1 FE_PHC2539_n1297 (.Y(FE_PHN2539_n1297), 
	.A(FE_PHN4014_n1297));
   DLY4X1 FE_PHC2538_n1824 (.Y(FE_PHN2538_n1824), 
	.A(FE_PHN3938_n1824));
   DLY4X1 FE_PHC2537_n2040 (.Y(FE_PHN2537_n2040), 
	.A(FE_PHN4172_n2040));
   DLY4X1 FE_PHC2536_n1809 (.Y(FE_PHN2536_n1809), 
	.A(n1809));
   DLY4X1 FE_PHC2535_n2239 (.Y(FE_PHN2535_n2239), 
	.A(FE_PHN4280_n2239));
   DLY4X1 FE_PHC2534_n2139 (.Y(FE_PHN2534_n2139), 
	.A(FE_PHN4603_n2139));
   DLY4X1 FE_PHC2533_n2148 (.Y(FE_PHN2533_n2148), 
	.A(FE_PHN4442_n2148));
   DLY4X1 FE_PHC2532_n1485 (.Y(FE_PHN2532_n1485), 
	.A(FE_PHN4104_n1485));
   DLY4X1 FE_PHC2531_n1460 (.Y(FE_PHN2531_n1460), 
	.A(n1460));
   DLY4X1 FE_PHC2530_n979 (.Y(FE_PHN2530_n979), 
	.A(FE_PHN4147_n979));
   DLY4X1 FE_PHC2529_n1695 (.Y(FE_PHN2529_n1695), 
	.A(FE_PHN4342_n1695));
   DLY4X1 FE_PHC2528_n1010 (.Y(FE_PHN2528_n1010), 
	.A(n1010));
   DLY4X1 FE_PHC2527_n1318 (.Y(FE_PHN2527_n1318), 
	.A(FE_PHN4090_n1318));
   DLY4X1 FE_PHC2526_n2049 (.Y(FE_PHN2526_n2049), 
	.A(FE_PHN4588_n2049));
   DLY4X1 FE_PHC2525_n1495 (.Y(FE_PHN2525_n1495), 
	.A(FE_PHN4013_n1495));
   DLY4X1 FE_PHC2524_n2254 (.Y(FE_PHN2524_n2254), 
	.A(FE_PHN3888_n2254));
   DLY4X1 FE_PHC2523_n1699 (.Y(FE_PHN2523_n1699), 
	.A(FE_PHN3925_n1699));
   DLY4X1 FE_PHC2522_n1900 (.Y(FE_PHN2522_n1900), 
	.A(FE_PHN4144_n1900));
   DLY4X1 FE_PHC2521_n2253 (.Y(FE_PHN2521_n2253), 
	.A(FE_PHN4331_n2253));
   DLY4X1 FE_PHC2520_n2191 (.Y(FE_PHN2520_n2191), 
	.A(FE_PHN4526_n2191));
   DLY4X1 FE_PHC2519_n2115 (.Y(FE_PHN2519_n2115), 
	.A(FE_PHN4267_n2115));
   DLY4X1 FE_PHC2518_n1310 (.Y(FE_PHN2518_n1310), 
	.A(FE_PHN3994_n1310));
   DLY4X1 FE_PHC2517_n941 (.Y(FE_PHN2517_n941), 
	.A(n941));
   DLY4X1 FE_PHC2516_n1761 (.Y(FE_PHN2516_n1761), 
	.A(n1761));
   DLY4X1 FE_PHC2515_n1740 (.Y(FE_PHN2515_n1740), 
	.A(FE_PHN4043_n1740));
   DLY4X1 FE_PHC2514_n1686 (.Y(FE_PHN2514_n1686), 
	.A(FE_PHN3987_n1686));
   DLY4X1 FE_PHC2513_n1903 (.Y(FE_PHN2513_n1903), 
	.A(FE_PHN4138_n1903));
   DLY4X1 FE_PHC2512_n922 (.Y(FE_PHN2512_n922), 
	.A(FE_PHN3942_n922));
   DLY4X1 FE_PHC2511_n1326 (.Y(FE_PHN2511_n1326), 
	.A(FE_PHN4799_n1326));
   DLY4X1 FE_PHC2510_n1274 (.Y(FE_PHN2510_n1274), 
	.A(FE_PHN4073_n1274));
   DLY4X1 FE_PHC2509_n976 (.Y(FE_PHN2509_n976), 
	.A(FE_PHN4294_n976));
   DLY4X1 FE_PHC2508_n2232 (.Y(FE_PHN2508_n2232), 
	.A(FE_PHN4435_n2232));
   DLY4X1 FE_PHC2507_n898 (.Y(FE_PHN2507_n898), 
	.A(FE_PHN3818_n898));
   DLY4X1 FE_PHC2506_n2123 (.Y(FE_PHN2506_n2123), 
	.A(FE_PHN4209_n2123));
   DLY4X1 FE_PHC2505_n1776 (.Y(FE_PHN2505_n1776), 
	.A(FE_PHN4378_n1776));
   DLY4X1 FE_PHC2504_n2174 (.Y(FE_PHN2504_n2174), 
	.A(FE_PHN4359_n2174));
   DLY4X1 FE_PHC2503_n897 (.Y(FE_PHN2503_n897), 
	.A(FE_PHN4015_n897));
   DLY4X1 FE_PHC2502_n2248 (.Y(FE_PHN2502_n2248), 
	.A(FE_PHN4101_n2248));
   DLY4X1 FE_PHC2501_n1731 (.Y(FE_PHN2501_n1731), 
	.A(FE_PHN4498_n1731));
   DLY4X1 FE_PHC2500_n2230 (.Y(FE_PHN2500_n2230), 
	.A(FE_PHN3882_n2230));
   DLY4X1 FE_PHC2499_n2277 (.Y(FE_PHN2499_n2277), 
	.A(n2277));
   DLY4X1 FE_PHC2498_n1861 (.Y(FE_PHN2498_n1861), 
	.A(FE_PHN4347_n1861));
   DLY4X1 FE_PHC2497_n1367 (.Y(FE_PHN2497_n1367), 
	.A(FE_PHN3993_n1367));
   DLY4X1 FE_PHC2496_n1670 (.Y(FE_PHN2496_n1670), 
	.A(FE_PHN4332_n1670));
   DLY4X1 FE_PHC2495_n980 (.Y(FE_PHN2495_n980), 
	.A(FE_PHN3845_n980));
   DLY4X1 FE_PHC2494_n1841 (.Y(FE_PHN2494_n1841), 
	.A(FE_PHN4205_n1841));
   DLY4X1 FE_PHC2493_n893 (.Y(FE_PHN2493_n893), 
	.A(FE_PHN3797_n893));
   DLY4X1 FE_PHC2492_n1478 (.Y(FE_PHN2492_n1478), 
	.A(FE_PHN4389_n1478));
   DLY4X1 FE_PHC2491_n1875 (.Y(FE_PHN2491_n1875), 
	.A(FE_PHN4000_n1875));
   DLY4X1 FE_PHC2490_n1884 (.Y(FE_PHN2490_n1884), 
	.A(FE_PHN4110_n1884));
   DLY4X1 FE_PHC2489_n921 (.Y(FE_PHN2489_n921), 
	.A(FE_PHN4404_n921));
   DLY4X1 FE_PHC2488_n2258 (.Y(FE_PHN2488_n2258), 
	.A(FE_PHN4297_n2258));
   DLY4X1 FE_PHC2487_n904 (.Y(FE_PHN2487_n904), 
	.A(FE_PHN4126_n904));
   DLY4X1 FE_PHC2486_n1842 (.Y(FE_PHN2486_n1842), 
	.A(FE_PHN3839_n1842));
   DLY4X1 FE_PHC2485_n1414 (.Y(FE_PHN2485_n1414), 
	.A(FE_PHN4340_n1414));
   DLY4X1 FE_PHC2484_n1725 (.Y(FE_PHN2484_n1725), 
	.A(FE_PHN4055_n1725));
   DLY4X1 FE_PHC2483_n1845 (.Y(FE_PHN2483_n1845), 
	.A(FE_PHN4290_n1845));
   DLY4X1 FE_PHC2482_n2072 (.Y(FE_PHN2482_n2072), 
	.A(FE_PHN3891_n2072));
   DLY4X1 FE_PHC2481_n996 (.Y(FE_PHN2481_n996), 
	.A(FE_PHN4041_n996));
   DLY4X1 FE_PHC2480_n912 (.Y(FE_PHN2480_n912), 
	.A(FE_PHN4496_n912));
   DLY4X1 FE_PHC2479_n982 (.Y(FE_PHN2479_n982), 
	.A(FE_PHN3976_n982));
   DLY4X1 FE_PHC2478_n1524 (.Y(FE_PHN2478_n1524), 
	.A(FE_PHN3924_n1524));
   DLY4X1 FE_PHC2477_n2037 (.Y(FE_PHN2477_n2037), 
	.A(n2037));
   DLY4X1 FE_PHC2476_n2208 (.Y(FE_PHN2476_n2208), 
	.A(FE_PHN3870_n2208));
   DLY4X1 FE_PHC2475_n951 (.Y(FE_PHN2475_n951), 
	.A(FE_PHN3957_n951));
   DLY4X1 FE_PHC2474_n1897 (.Y(FE_PHN2474_n1897), 
	.A(n1897));
   DLY4X1 FE_PHC2473_n1747 (.Y(FE_PHN2473_n1747), 
	.A(FE_PHN3937_n1747));
   DLY4X1 FE_PHC2472_n2150 (.Y(FE_PHN2472_n2150), 
	.A(FE_PHN3802_n2150));
   DLY4X1 FE_PHC2471_n2209 (.Y(FE_PHN2471_n2209), 
	.A(FE_PHN4718_n2209));
   DLY4X1 FE_PHC2470_n2118 (.Y(FE_PHN2470_n2118), 
	.A(FE_PHN3899_n2118));
   DLY4X1 FE_PHC2469_n1314 (.Y(FE_PHN2469_n1314), 
	.A(FE_PHN4019_n1314));
   DLY4X1 FE_PHC2468_n952 (.Y(FE_PHN2468_n952), 
	.A(FE_PHN4233_n952));
   DLY4X1 FE_PHC2467_n1795 (.Y(FE_PHN2467_n1795), 
	.A(FE_PHN3940_n1795));
   DLY4X1 FE_PHC2466_n2262 (.Y(FE_PHN2466_n2262), 
	.A(FE_PHN3988_n2262));
   DLY4X1 FE_PHC2465_n924 (.Y(FE_PHN2465_n924), 
	.A(n924));
   DLY4X1 FE_PHC2464_n1701 (.Y(FE_PHN2464_n1701), 
	.A(FE_PHN3887_n1701));
   DLY4X1 FE_PHC2463_n1404 (.Y(FE_PHN2463_n1404), 
	.A(FE_PHN3773_n1404));
   DLY4X1 FE_PHC2462_n1857 (.Y(FE_PHN2462_n1857), 
	.A(FE_PHN4580_n1857));
   DLY4X1 FE_PHC2461_n1882 (.Y(FE_PHN2461_n1882), 
	.A(FE_PHN3766_n1882));
   DLY4X1 FE_PHC2460_n1000 (.Y(FE_PHN2460_n1000), 
	.A(FE_PHN3939_n1000));
   DLY4X1 FE_PHC2459_n1006 (.Y(FE_PHN2459_n1006), 
	.A(FE_PHN4543_n1006));
   DLY4X1 FE_PHC2458_n1334 (.Y(FE_PHN2458_n1334), 
	.A(FE_PHN4068_n1334));
   DLY4X1 FE_PHC2457_n889 (.Y(FE_PHN2457_n889), 
	.A(FE_PHN3877_n889));
   DLY4X1 FE_PHC2456_n2173 (.Y(FE_PHN2456_n2173), 
	.A(FE_PHN3860_n2173));
   DLY4X1 FE_PHC2455_n2275 (.Y(FE_PHN2455_n2275), 
	.A(FE_PHN4631_n2275));
   DLY4X1 FE_PHC2454_n1680 (.Y(FE_PHN2454_n1680), 
	.A(FE_PHN3970_n1680));
   DLY4X1 FE_PHC2453_n2103 (.Y(FE_PHN2453_n2103), 
	.A(FE_PHN3886_n2103));
   DLY4X1 FE_PHC2452_n2162 (.Y(FE_PHN2452_n2162), 
	.A(FE_PHN4005_n2162));
   DLY4X1 FE_PHC2451_n1806 (.Y(FE_PHN2451_n1806), 
	.A(FE_PHN4622_n1806));
   DLY4X1 FE_PHC2450_n1772 (.Y(FE_PHN2450_n1772), 
	.A(FE_PHN3962_n1772));
   DLY4X1 FE_PHC2449_n2135 (.Y(FE_PHN2449_n2135), 
	.A(FE_PHN4009_n2135));
   DLY4X1 FE_PHC2448_n1698 (.Y(FE_PHN2448_n1698), 
	.A(FE_PHN3971_n1698));
   DLY4X1 FE_PHC2447_n1892 (.Y(FE_PHN2447_n1892), 
	.A(FE_PHN4385_n1892));
   DLY4X1 FE_PHC2446_n1401 (.Y(FE_PHN2446_n1401), 
	.A(FE_PHN4434_n1401));
   DLY4X1 FE_PHC2445_n1328 (.Y(FE_PHN2445_n1328), 
	.A(FE_PHN3723_n1328));
   DLY4X1 FE_PHC2444_n1433 (.Y(FE_PHN2444_n1433), 
	.A(FE_PHN3966_n1433));
   DLY4X1 FE_PHC2443_n2108 (.Y(FE_PHN2443_n2108), 
	.A(FE_PHN3959_n2108));
   DLY4X1 FE_PHC2442_n1681 (.Y(FE_PHN2442_n1681), 
	.A(FE_PHN4807_n1681));
   DLY4X1 FE_PHC2441_n1434 (.Y(FE_PHN2441_n1434), 
	.A(n1434));
   DLY4X1 FE_PHC2440_n901 (.Y(FE_PHN2440_n901), 
	.A(n901));
   DLY4X1 FE_PHC2439_n2207 (.Y(FE_PHN2439_n2207), 
	.A(FE_PHN4257_n2207));
   DLY4X1 FE_PHC2438_n1822 (.Y(FE_PHN2438_n1822), 
	.A(FE_PHN3812_n1822));
   DLY4X1 FE_PHC2437_n1723 (.Y(FE_PHN2437_n1723), 
	.A(FE_PHN3799_n1723));
   DLY4X1 FE_PHC2436_n1735 (.Y(FE_PHN2436_n1735), 
	.A(FE_PHN4223_n1735));
   DLY4X1 FE_PHC2435_n1797 (.Y(FE_PHN2435_n1797), 
	.A(FE_PHN3896_n1797));
   DLY4X1 FE_PHC2434_n969 (.Y(FE_PHN2434_n969), 
	.A(FE_PHN4798_n969));
   DLY4X1 FE_PHC2433_n966 (.Y(FE_PHN2433_n966), 
	.A(FE_PHN4046_n966));
   DLY4X1 FE_PHC2432_n1780 (.Y(FE_PHN2432_n1780), 
	.A(FE_PHN4221_n1780));
   DLY4X1 FE_PHC2431_n950 (.Y(FE_PHN2431_n950), 
	.A(FE_PHN4039_n950));
   DLY4X1 FE_PHC2430_n1673 (.Y(FE_PHN2430_n1673), 
	.A(FE_PHN3805_n1673));
   DLY4X1 FE_PHC2429_n1821 (.Y(FE_PHN2429_n1821), 
	.A(FE_PHN3945_n1821));
   DLY4X1 FE_PHC2428_n1858 (.Y(FE_PHN2428_n1858), 
	.A(FE_PHN3913_n1858));
   DLY4X1 FE_PHC2427_n2051 (.Y(FE_PHN2427_n2051), 
	.A(FE_PHN3895_n2051));
   DLY4X1 FE_PHC2426_n1697 (.Y(FE_PHN2426_n1697), 
	.A(FE_PHN4353_n1697));
   DLY4X1 FE_PHC2425_n1748 (.Y(FE_PHN2425_n1748), 
	.A(FE_PHN4249_n1748));
   DLY4X1 FE_PHC2424_n2159 (.Y(FE_PHN2424_n2159), 
	.A(FE_PHN4487_n2159));
   DLY4X1 FE_PHC2423_n1707 (.Y(FE_PHN2423_n1707), 
	.A(FE_PHN4224_n1707));
   DLY4X1 FE_PHC2422_n1702 (.Y(FE_PHN2422_n1702), 
	.A(FE_PHN3904_n1702));
   DLY4X1 FE_PHC2421_n1831 (.Y(FE_PHN2421_n1831), 
	.A(FE_PHN4177_n1831));
   DLY4X1 FE_PHC2420_n1683 (.Y(FE_PHN2420_n1683), 
	.A(FE_PHN4451_n1683));
   DLY4X1 FE_PHC2419_n1830 (.Y(FE_PHN2419_n1830), 
	.A(FE_PHN4218_n1830));
   DLY4X1 FE_PHC2418_n938 (.Y(FE_PHN2418_n938), 
	.A(FE_PHN3880_n938));
   DLY4X1 FE_PHC2417_n895 (.Y(FE_PHN2417_n895), 
	.A(FE_PHN4124_n895));
   DLY4X1 FE_PHC2416_n1519 (.Y(FE_PHN2416_n1519), 
	.A(FE_PHN4056_n1519));
   DLY4X1 FE_PHC2415_n2276 (.Y(FE_PHN2415_n2276), 
	.A(FE_PHN3785_n2276));
   DLY4X1 FE_PHC2414_n1869 (.Y(FE_PHN2414_n1869), 
	.A(FE_PHN3926_n1869));
   DLY4X1 FE_PHC2413_n1837 (.Y(FE_PHN2413_n1837), 
	.A(FE_PHN4199_n1837));
   DLY4X1 FE_PHC2412_n2236 (.Y(FE_PHN2412_n2236), 
	.A(FE_PHN4081_n2236));
   DLY4X1 FE_PHC2411_n906 (.Y(FE_PHN2411_n906), 
	.A(n906));
   DLY4X1 FE_PHC2410_n2043 (.Y(FE_PHN2410_n2043), 
	.A(FE_PHN4163_n2043));
   DLY4X1 FE_PHC2409_n1815 (.Y(FE_PHN2409_n1815), 
	.A(FE_PHN3946_n1815));
   DLY4X1 FE_PHC2408_n2184 (.Y(FE_PHN2408_n2184), 
	.A(FE_PHN4254_n2184));
   DLY4X1 FE_PHC2407_n1448 (.Y(FE_PHN2407_n1448), 
	.A(FE_PHN3897_n1448));
   DLY4X1 FE_PHC2406_n2161 (.Y(FE_PHN2406_n2161), 
	.A(n2161));
   DLY4X1 FE_PHC2405_n964 (.Y(FE_PHN2405_n964), 
	.A(FE_PHN3853_n964));
   DLY4X1 FE_PHC2404_n1513 (.Y(FE_PHN2404_n1513), 
	.A(FE_PHN4089_n1513));
   DLY4X1 FE_PHC2403_n2087 (.Y(FE_PHN2403_n2087), 
	.A(FE_PHN3923_n2087));
   DLY4X1 FE_PHC2402_n1743 (.Y(FE_PHN2402_n1743), 
	.A(FE_PHN3862_n1743));
   DLY4X1 FE_PHC2401_n1398 (.Y(FE_PHN2401_n1398), 
	.A(n1398));
   DLY4X1 FE_PHC2400_n1003 (.Y(FE_PHN2400_n1003), 
	.A(n1003));
   DLY4X1 FE_PHC2399_n1484 (.Y(FE_PHN2399_n1484), 
	.A(FE_PHN4251_n1484));
   DLY4X1 FE_PHC2398_n1781 (.Y(FE_PHN2398_n1781), 
	.A(FE_PHN3808_n1781));
   DLY4X1 FE_PHC2397_n1783 (.Y(FE_PHN2397_n1783), 
	.A(FE_PHN4230_n1783));
   DLY4X1 FE_PHC2396_n1654 (.Y(FE_PHN2396_n1654), 
	.A(FE_PHN4283_n1654));
   DLY4X1 FE_PHC2395_n1483 (.Y(FE_PHN2395_n1483), 
	.A(FE_PHN3984_n1483));
   DLY4X1 FE_PHC2394_n1865 (.Y(FE_PHN2394_n1865), 
	.A(FE_PHN4475_n1865));
   DLY4X1 FE_PHC2393_n890 (.Y(FE_PHN2393_n890), 
	.A(FE_PHN4048_n890));
   DLY4X1 FE_PHC2392_n2153 (.Y(FE_PHN2392_n2153), 
	.A(FE_PHN4120_n2153));
   DLY4X1 FE_PHC2391_n1472 (.Y(FE_PHN2391_n1472), 
	.A(FE_PHN3868_n1472));
   DLY4X1 FE_PHC2390_n2134 (.Y(FE_PHN2390_n2134), 
	.A(FE_PHN3741_n2134));
   DLY4X1 FE_PHC2389_n1410 (.Y(FE_PHN2389_n1410), 
	.A(FE_PHN4141_n1410));
   DLY4X1 FE_PHC2388_n2216 (.Y(FE_PHN2388_n2216), 
	.A(FE_PHN4133_n2216));
   DLY4X1 FE_PHC2387_n2194 (.Y(FE_PHN2387_n2194), 
	.A(FE_PHN4384_n2194));
   DLY4X1 FE_PHC2386_n2269 (.Y(FE_PHN2386_n2269), 
	.A(FE_PHN3809_n2269));
   DLY4X1 FE_PHC2385_n1709 (.Y(FE_PHN2385_n1709), 
	.A(FE_PHN3955_n1709));
   DLY4X1 FE_PHC2384_n1474 (.Y(FE_PHN2384_n1474), 
	.A(FE_PHN4008_n1474));
   DLY4X1 FE_PHC2383_n1711 (.Y(FE_PHN2383_n1711), 
	.A(FE_PHN3901_n1711));
   DLY4X1 FE_PHC2382_n1870 (.Y(FE_PHN2382_n1870), 
	.A(FE_PHN3826_n1870));
   DLY4X1 FE_PHC2381_n2167 (.Y(FE_PHN2381_n2167), 
	.A(FE_PHN4450_n2167));
   DLY4X1 FE_PHC2380_n1458 (.Y(FE_PHN2380_n1458), 
	.A(FE_PHN3749_n1458));
   DLY4X1 FE_PHC2379_n2233 (.Y(FE_PHN2379_n2233), 
	.A(FE_PHN3843_n2233));
   DLY4X1 FE_PHC2378_n1466 (.Y(FE_PHN2378_n1466), 
	.A(FE_PHN4037_n1466));
   DLY4X1 FE_PHC2377_n2085 (.Y(FE_PHN2377_n2085), 
	.A(FE_PHN4050_n2085));
   DLY4X1 FE_PHC2376_n1502 (.Y(FE_PHN2376_n1502), 
	.A(FE_PHN3801_n1502));
   DLY4X1 FE_PHC2375_n1881 (.Y(FE_PHN2375_n1881), 
	.A(FE_PHN4250_n1881));
   DLY4X1 FE_PHC2374_n2226 (.Y(FE_PHN2374_n2226), 
	.A(FE_PHN4266_n2226));
   DLY4X1 FE_PHC2373_n1798 (.Y(FE_PHN2373_n1798), 
	.A(FE_PHN3752_n1798));
   DLY4X1 FE_PHC2372_n2075 (.Y(FE_PHN2372_n2075), 
	.A(FE_PHN3832_n2075));
   DLY4X1 FE_PHC2371_n1819 (.Y(FE_PHN2371_n1819), 
	.A(n1819));
   DLY4X1 FE_PHC2370_n1694 (.Y(FE_PHN2370_n1694), 
	.A(FE_PHN3706_n1694));
   DLY4X1 FE_PHC2369_n1828 (.Y(FE_PHN2369_n1828), 
	.A(FE_PHN4188_n1828));
   DLY4X1 FE_PHC2368_n1899 (.Y(FE_PHN2368_n1899), 
	.A(FE_PHN4069_n1899));
   DLY4X1 FE_PHC2367_n2222 (.Y(FE_PHN2367_n2222), 
	.A(FE_PHN4158_n2222));
   DLY4X1 FE_PHC2366_n1755 (.Y(FE_PHN2366_n1755), 
	.A(FE_PHN4502_n1755));
   DLY4X1 FE_PHC2365_n1741 (.Y(FE_PHN2365_n1741), 
	.A(FE_PHN4026_n1741));
   DLY4X1 FE_PHC2364_n1421 (.Y(FE_PHN2364_n1421), 
	.A(n1421));
   DLY4X1 FE_PHC2363_n2245 (.Y(FE_PHN2363_n2245), 
	.A(FE_PHN3849_n2245));
   DLY4X1 FE_PHC2362_n1465 (.Y(FE_PHN2362_n1465), 
	.A(FE_PHN3767_n1465));
   DLY4X1 FE_PHC2361_n2071 (.Y(FE_PHN2361_n2071), 
	.A(FE_PHN4202_n2071));
   DLY4X1 FE_PHC2360_n1742 (.Y(FE_PHN2360_n1742), 
	.A(FE_PHN4162_n1742));
   DLY4X1 FE_PHC2359_n2080 (.Y(FE_PHN2359_n2080), 
	.A(FE_PHN3804_n2080));
   DLY4X1 FE_PHC2358_n1523 (.Y(FE_PHN2358_n1523), 
	.A(FE_PHN3840_n1523));
   DLY4X1 FE_PHC2357_n2278 (.Y(FE_PHN2357_n2278), 
	.A(FE_PHN4179_n2278));
   DLY4X1 FE_PHC2356_n1504 (.Y(FE_PHN2356_n1504), 
	.A(FE_PHN4178_n1504));
   DLY4X1 FE_PHC2355_n2127 (.Y(FE_PHN2355_n2127), 
	.A(FE_PHN3985_n2127));
   DLY4X1 FE_PHC2354_n2130 (.Y(FE_PHN2354_n2130), 
	.A(FE_PHN3806_n2130));
   DLY4X1 FE_PHC2353_n1437 (.Y(FE_PHN2353_n1437), 
	.A(FE_PHN3833_n1437));
   DLY4X1 FE_PHC2352_n2227 (.Y(FE_PHN2352_n2227), 
	.A(FE_PHN3751_n2227));
   DLY4X1 FE_PHC2351_n2252 (.Y(FE_PHN2351_n2252), 
	.A(FE_PHN3997_n2252));
   DLY4X1 FE_PHC2350_n1674 (.Y(FE_PHN2350_n1674), 
	.A(n1674));
   DLY4X1 FE_PHC2349_n1457 (.Y(FE_PHN2349_n1457), 
	.A(FE_PHN4112_n1457));
   DLY4X1 FE_PHC2348_n1719 (.Y(FE_PHN2348_n1719), 
	.A(FE_PHN3793_n1719));
   DLY4X1 FE_PHC2347_n2041 (.Y(FE_PHN2347_n2041), 
	.A(FE_PHN3914_n2041));
   DLY4X1 FE_PHC2346_n2270 (.Y(FE_PHN2346_n2270), 
	.A(FE_PHN3873_n2270));
   DLY4X1 FE_PHC2345_n2203 (.Y(FE_PHN2345_n2203), 
	.A(FE_PHN3828_n2203));
   DLY4X1 FE_PHC2344_n2113 (.Y(FE_PHN2344_n2113), 
	.A(FE_PHN3673_n2113));
   DLY4X1 FE_PHC2343_n1883 (.Y(FE_PHN2343_n1883), 
	.A(FE_PHN3905_n1883));
   DLY4X1 FE_PHC2342_n2128 (.Y(FE_PHN2342_n2128), 
	.A(FE_PHN4099_n2128));
   DLY4X1 FE_PHC2341_n2052 (.Y(FE_PHN2341_n2052), 
	.A(FE_PHN4193_n2052));
   DLY4X1 FE_PHC2340_n2102 (.Y(FE_PHN2340_n2102), 
	.A(FE_PHN4011_n2102));
   DLY4X1 FE_PHC2339_n2112 (.Y(FE_PHN2339_n2112), 
	.A(FE_PHN3712_n2112));
   DLY4X1 FE_PHC2338_n1893 (.Y(FE_PHN2338_n1893), 
	.A(FE_PHN3683_n1893));
   DLY4X1 FE_PHC2337_n1791 (.Y(FE_PHN2337_n1791), 
	.A(FE_PHN4330_n1791));
   DLY4X1 FE_PHC2336_n1794 (.Y(FE_PHN2336_n1794), 
	.A(FE_PHN3675_n1794));
   DLY4X1 FE_PHC2335_n1777 (.Y(FE_PHN2335_n1777), 
	.A(FE_PHN4109_n1777));
   DLY4X1 FE_PHC2334_n2156 (.Y(FE_PHN2334_n2156), 
	.A(FE_PHN4279_n2156));
   DLY4X1 FE_PHC2333_n2217 (.Y(FE_PHN2333_n2217), 
	.A(FE_PHN3714_n2217));
   DLY4X1 FE_PHC2332_n1811 (.Y(FE_PHN2332_n1811), 
	.A(n1811));
   DLY4X1 FE_PHC2331_n1726 (.Y(FE_PHN2331_n1726), 
	.A(FE_PHN3779_n1726));
   DLY4X1 FE_PHC2330_n1778 (.Y(FE_PHN2330_n1778), 
	.A(FE_PHN3872_n1778));
   DLY4X1 FE_PHC2329_n2225 (.Y(FE_PHN2329_n2225), 
	.A(FE_PHN3852_n2225));
   DLY4X1 FE_PHC2328_n2213 (.Y(FE_PHN2328_n2213), 
	.A(FE_PHN3780_n2213));
   DLY4X1 FE_PHC2327_n1453 (.Y(FE_PHN2327_n1453), 
	.A(n1453));
   DLY4X1 FE_PHC2326_n1514 (.Y(FE_PHN2326_n1514), 
	.A(FE_PHN4461_n1514));
   DLY4X1 FE_PHC2325_n2110 (.Y(FE_PHN2325_n2110), 
	.A(FE_PHN3972_n2110));
   DLY4X1 FE_PHC2324_n2053 (.Y(FE_PHN2324_n2053), 
	.A(n2053));
   DLY4X1 FE_PHC2323_n1411 (.Y(FE_PHN2323_n1411), 
	.A(FE_PHN3747_n1411));
   DLY4X1 FE_PHC2322_n1512 (.Y(FE_PHN2322_n1512), 
	.A(FE_PHN3709_n1512));
   DLY4X1 FE_PHC2321_n1851 (.Y(FE_PHN2321_n1851), 
	.A(FE_PHN4121_n1851));
   DLY4X1 FE_PHC2320_n1901 (.Y(FE_PHN2320_n1901), 
	.A(n1901));
   DLY4X1 FE_PHC2319_n2268 (.Y(FE_PHN2319_n2268), 
	.A(FE_PHN3990_n2268));
   DLY4X1 FE_PHC2318_n1767 (.Y(FE_PHN2318_n1767), 
	.A(FE_PHN4376_n1767));
   DLY4X1 FE_PHC2317_n1507 (.Y(FE_PHN2317_n1507), 
	.A(FE_PHN4171_n1507));
   DLY4X1 FE_PHC2316_n2244 (.Y(FE_PHN2316_n2244), 
	.A(FE_PHN3874_n2244));
   DLY4X1 FE_PHC2315_n1860 (.Y(FE_PHN2315_n1860), 
	.A(FE_PHN3770_n1860));
   DLY4X1 FE_PHC2314_n1684 (.Y(FE_PHN2314_n1684), 
	.A(FE_PHN3918_n1684));
   DLY4X1 FE_PHC2313_n1677 (.Y(FE_PHN2313_n1677), 
	.A(FE_PHN4148_n1677));
   DLY4X1 FE_PHC2312_n1475 (.Y(FE_PHN2312_n1475), 
	.A(n1475));
   DLY4X1 FE_PHC2311_n1757 (.Y(FE_PHN2311_n1757), 
	.A(FE_PHN4030_n1757));
   DLY4X1 FE_PHC2310_n2177 (.Y(FE_PHN2310_n2177), 
	.A(FE_PHN3831_n2177));
   DLY4X1 FE_PHC2309_n1854 (.Y(FE_PHN2309_n1854), 
	.A(FE_PHN4023_n1854));
   DLY4X1 FE_PHC2308_n2086 (.Y(FE_PHN2308_n2086), 
	.A(FE_PHN3796_n2086));
   DLY4X1 FE_PHC2307_n2257 (.Y(FE_PHN2307_n2257), 
	.A(FE_PHN3995_n2257));
   DLY4X1 FE_PHC2306_n1728 (.Y(FE_PHN2306_n1728), 
	.A(FE_PHN4513_n1728));
   DLY4X1 FE_PHC2305_n1480 (.Y(FE_PHN2305_n1480), 
	.A(FE_PHN4232_n1480));
   DLY4X1 FE_PHC2304_n2292 (.Y(FE_PHN2304_n2292), 
	.A(FE_PHN4078_n2292));
   DLY4X1 FE_PHC2303_n1906 (.Y(FE_PHN2303_n1906), 
	.A(FE_PHN3810_n1906));
   DLY4X1 FE_PHC2302_n1436 (.Y(FE_PHN2302_n1436), 
	.A(FE_PHN3721_n1436));
   DLY4X1 FE_PHC2301_n2078 (.Y(FE_PHN2301_n2078), 
	.A(FE_PHN3745_n2078));
   DLY4X1 FE_PHC2300_n1469 (.Y(FE_PHN2300_n1469), 
	.A(FE_PHN4113_n1469));
   DLY4X1 FE_PHC2299_n1488 (.Y(FE_PHN2299_n1488), 
	.A(FE_PHN4808_n1488));
   DLY4X1 FE_PHC2298_n1409 (.Y(FE_PHN2298_n1409), 
	.A(FE_PHN4161_n1409));
   DLY4X1 FE_PHC2297_n1415 (.Y(FE_PHN2297_n1415), 
	.A(FE_PHN3820_n1415));
   DLY4X1 FE_PHC2296_n1441 (.Y(FE_PHN2296_n1441), 
	.A(FE_PHN3920_n1441));
   DLY4X1 FE_PHC2295_n1672 (.Y(FE_PHN2295_n1672), 
	.A(FE_PHN3813_n1672));
   DLY4X1 FE_PHC2294_n2074 (.Y(FE_PHN2294_n2074), 
	.A(FE_PHN3715_n2074));
   DLY4X1 FE_PHC2293_n2095 (.Y(FE_PHN2293_n2095), 
	.A(FE_PHN3982_n2095));
   DLY4X1 FE_PHC2292_n2238 (.Y(FE_PHN2292_n2238), 
	.A(FE_PHN4479_n2238));
   DLY4X1 FE_PHC2291_n1664 (.Y(FE_PHN2291_n1664), 
	.A(FE_PHN3968_n1664));
   DLY4X1 FE_PHC2290_n1454 (.Y(FE_PHN2290_n1454), 
	.A(FE_PHN3679_n1454));
   DLY4X1 FE_PHC2289_n1473 (.Y(FE_PHN2289_n1473), 
	.A(FE_PHN3803_n1473));
   DLY4X1 FE_PHC2288_n1399 (.Y(FE_PHN2288_n1399), 
	.A(FE_PHN3788_n1399));
   DLY4X1 FE_PHC2287_n2155 (.Y(FE_PHN2287_n2155), 
	.A(FE_PHN4616_n2155));
   DLY4X1 FE_PHC2286_n2272 (.Y(FE_PHN2286_n2272), 
	.A(FE_PHN3943_n2272));
   DLY4X1 FE_PHC2285_n1429 (.Y(FE_PHN2285_n1429), 
	.A(FE_PHN3718_n1429));
   DLY4X1 FE_PHC2284_n1876 (.Y(FE_PHN2284_n1876), 
	.A(FE_PHN3912_n1876));
   DLY4X1 FE_PHC2283_n2164 (.Y(FE_PHN2283_n2164), 
	.A(FE_PHN4106_n2164));
   DLY4X1 FE_PHC2282_n1770 (.Y(FE_PHN2282_n1770), 
	.A(FE_PHN4071_n1770));
   DLY4X1 FE_PHC2281_n1462 (.Y(FE_PHN2281_n1462), 
	.A(FE_PHN4529_n1462));
   DLY4X1 FE_PHC2280_n2101 (.Y(FE_PHN2280_n2101), 
	.A(FE_PHN4033_n2101));
   DLY4X1 FE_PHC2279_n2202 (.Y(FE_PHN2279_n2202), 
	.A(FE_PHN3783_n2202));
   DLY4X1 FE_PHC2278_n2145 (.Y(FE_PHN2278_n2145), 
	.A(FE_PHN3725_n2145));
   DLY4X1 FE_PHC2277_n1907 (.Y(FE_PHN2277_n1907), 
	.A(FE_PHN4131_n1907));
   DLY4X1 FE_PHC2276_n2093 (.Y(FE_PHN2276_n2093), 
	.A(FE_PHN4169_n2093));
   DLY4X1 FE_PHC2275_n2186 (.Y(FE_PHN2275_n2186), 
	.A(n2186));
   DLY4X1 FE_PHC2274_n1508 (.Y(FE_PHN2274_n1508), 
	.A(FE_PHN3771_n1508));
   DLY4X1 FE_PHC2273_n1506 (.Y(FE_PHN2273_n1506), 
	.A(FE_PHN3859_n1506));
   DLY4X1 FE_PHC2272_n1467 (.Y(FE_PHN2272_n1467), 
	.A(FE_PHN3989_n1467));
   DLY4X1 FE_PHC2271_n1890 (.Y(FE_PHN2271_n1890), 
	.A(FE_PHN3998_n1890));
   DLY4X1 FE_PHC2270_n1682 (.Y(FE_PHN2270_n1682), 
	.A(FE_PHN3649_n1682));
   DLY4X1 FE_PHC2269_n2283 (.Y(FE_PHN2269_n2283), 
	.A(FE_PHN4608_n2283));
   DLY4X1 FE_PHC2268_n1662 (.Y(FE_PHN2268_n1662), 
	.A(FE_PHN3816_n1662));
   DLY4X1 FE_PHC2267_n1721 (.Y(FE_PHN2267_n1721), 
	.A(FE_PHN3719_n1721));
   DLY4X1 FE_PHC2266_n1823 (.Y(FE_PHN2266_n1823), 
	.A(FE_PHN3726_n1823));
   DLY4X1 FE_PHC2265_n1521 (.Y(FE_PHN2265_n1521), 
	.A(FE_PHN3950_n1521));
   DLY4X1 FE_PHC2264_n1503 (.Y(FE_PHN2264_n1503), 
	.A(FE_PHN3660_n1503));
   DLY4X1 FE_PHC2263_n1463 (.Y(FE_PHN2263_n1463), 
	.A(FE_PHN3684_n1463));
   DLY4X1 FE_PHC2262_n1443 (.Y(FE_PHN2262_n1443), 
	.A(FE_PHN3756_n1443));
   DLY4X1 FE_PHC2261_n2140 (.Y(FE_PHN2261_n2140), 
	.A(FE_PHN4259_n2140));
   DLY4X1 FE_PHC2260_n2201 (.Y(FE_PHN2260_n2201), 
	.A(FE_PHN4692_n2201));
   DLY4X1 FE_PHC2259_n1665 (.Y(FE_PHN2259_n1665), 
	.A(FE_PHN4132_n1665));
   DLY4X1 FE_PHC2258_n2240 (.Y(FE_PHN2258_n2240), 
	.A(FE_PHN4077_n2240));
   DLY4X1 FE_PHC2257_n2247 (.Y(FE_PHN2257_n2247), 
	.A(FE_PHN3655_n2247));
   DLY4X1 FE_PHC2256_n1801 (.Y(FE_PHN2256_n1801), 
	.A(FE_PHN3750_n1801));
   DLY4X1 FE_PHC2255_n1693 (.Y(FE_PHN2255_n1693), 
	.A(FE_PHN3659_n1693));
   DLY4X1 FE_PHC2254_n2100 (.Y(FE_PHN2254_n2100), 
	.A(FE_PHN4029_n2100));
   DLY4X1 FE_PHC2253_n2192 (.Y(FE_PHN2253_n2192), 
	.A(FE_PHN3944_n2192));
   DLY4X1 FE_PHC2252_n1756 (.Y(FE_PHN2252_n1756), 
	.A(FE_PHN3772_n1756));
   DLY4X1 FE_PHC2251_n2067 (.Y(FE_PHN2251_n2067), 
	.A(FE_PHN3823_n2067));
   DLY4X1 FE_PHC2250_n1862 (.Y(FE_PHN2250_n1862), 
	.A(FE_PHN4076_n1862));
   DLY4X1 FE_PHC2249_n1779 (.Y(FE_PHN2249_n1779), 
	.A(FE_PHN4476_n1779));
   DLY4X1 FE_PHC2248_n2131 (.Y(FE_PHN2248_n2131), 
	.A(FE_PHN4130_n2131));
   DLY4X1 FE_PHC2247_n2083 (.Y(FE_PHN2247_n2083), 
	.A(FE_PHN3764_n2083));
   DLY4X1 FE_PHC2246_n1685 (.Y(FE_PHN2246_n1685), 
	.A(FE_PHN3667_n1685));
   DLY4X1 FE_PHC2245_n2090 (.Y(FE_PHN2245_n2090), 
	.A(FE_PHN4063_n2090));
   DLY4X1 FE_PHC2244_n2097 (.Y(FE_PHN2244_n2097), 
	.A(FE_PHN3777_n2097));
   DLY4X1 FE_PHC2243_n1866 (.Y(FE_PHN2243_n1866), 
	.A(FE_PHN4036_n1866));
   DLY4X1 FE_PHC2242_n1817 (.Y(FE_PHN2242_n1817), 
	.A(FE_PHN3790_n1817));
   DLY4X1 FE_PHC2241_n2220 (.Y(FE_PHN2241_n2220), 
	.A(FE_PHN3636_n2220));
   DLY4X1 FE_PHC2240_n1792 (.Y(FE_PHN2240_n1792), 
	.A(FE_PHN4070_n1792));
   DLY4X1 FE_PHC2239_n2055 (.Y(FE_PHN2239_n2055), 
	.A(FE_PHN3762_n2055));
   DLY4X1 FE_PHC2238_n1720 (.Y(FE_PHN2238_n1720), 
	.A(FE_PHN3630_n1720));
   DLY4X1 FE_PHC2237_n1509 (.Y(FE_PHN2237_n1509), 
	.A(FE_PHN3775_n1509));
   DLY4X1 FE_PHC2236_n1787 (.Y(FE_PHN2236_n1787), 
	.A(FE_PHN3748_n1787));
   DLY4X1 FE_PHC2235_n1727 (.Y(FE_PHN2235_n1727), 
	.A(FE_PHN3781_n1727));
   DLY4X1 FE_PHC2234_n1889 (.Y(FE_PHN2234_n1889), 
	.A(n1889));
   DLY4X1 FE_PHC2233_n1788 (.Y(FE_PHN2233_n1788), 
	.A(FE_PHN4105_n1788));
   DLY4X1 FE_PHC2232_n1785 (.Y(FE_PHN2232_n1785), 
	.A(n1785));
   DLY4X1 FE_PHC2231_n2165 (.Y(FE_PHN2231_n2165), 
	.A(n2165));
   DLY4X1 FE_PHC2230_n1868 (.Y(FE_PHN2230_n1868), 
	.A(FE_PHN3952_n1868));
   DLY4X1 FE_PHC2229_n1877 (.Y(FE_PHN2229_n1877), 
	.A(FE_PHN3906_n1877));
   DLY4X1 FE_PHC2228_n1451 (.Y(FE_PHN2228_n1451), 
	.A(FE_PHN3742_n1451));
   DLY4X1 FE_PHC2227_n2126 (.Y(FE_PHN2227_n2126), 
	.A(FE_PHN3635_n2126));
   DLY4X1 FE_PHC2226_n2224 (.Y(FE_PHN2226_n2224), 
	.A(FE_PHN3704_n2224));
   DLY4X1 FE_PHC2225_n2255 (.Y(FE_PHN2225_n2255), 
	.A(FE_PHN3627_n2255));
   DLY4X1 FE_PHC2224_n1456 (.Y(FE_PHN2224_n1456), 
	.A(FE_PHN4017_n1456));
   DLY4X1 FE_PHC2223_n1494 (.Y(FE_PHN2223_n1494), 
	.A(FE_PHN3759_n1494));
   DLY4X1 FE_PHC2222_n2274 (.Y(FE_PHN2222_n2274), 
	.A(n2274));
   DLY4X1 FE_PHC2221_n1803 (.Y(FE_PHN2221_n1803), 
	.A(FE_PHN3744_n1803));
   DLY4X1 FE_PHC2220_n2219 (.Y(FE_PHN2220_n2219), 
	.A(n2219));
   DLY4X1 FE_PHC2219_n1754 (.Y(FE_PHN2219_n1754), 
	.A(FE_PHN3757_n1754));
   DLY4X1 FE_PHC2218_n1898 (.Y(FE_PHN2218_n1898), 
	.A(FE_PHN3800_n1898));
   DLY4X1 FE_PHC2217_n2154 (.Y(FE_PHN2217_n2154), 
	.A(FE_PHN3637_n2154));
   DLY4X1 FE_PHC2216_n2250 (.Y(FE_PHN2216_n2250), 
	.A(FE_PHN3695_n2250));
   DLY4X1 FE_PHC2215_n2260 (.Y(FE_PHN2215_n2260), 
	.A(FE_PHN3732_n2260));
   DLY4X1 FE_PHC2214_n1863 (.Y(FE_PHN2214_n1863), 
	.A(FE_PHN3738_n1863));
   DLY4X1 FE_PHC2213_n1696 (.Y(FE_PHN2213_n1696), 
	.A(FE_PHN3969_n1696));
   DLY4X1 FE_PHC2212_n1844 (.Y(FE_PHN2212_n1844), 
	.A(FE_PHN3983_n1844));
   DLY4X1 FE_PHC2211_n2178 (.Y(FE_PHN2211_n2178), 
	.A(FE_PHN3746_n2178));
   DLY4X1 FE_PHC2210_n1832 (.Y(FE_PHN2210_n1832), 
	.A(FE_PHN4440_n1832));
   DLY4X1 FE_PHC2209_n2231 (.Y(FE_PHN2209_n2231), 
	.A(FE_PHN3632_n2231));
   DLY4X1 FE_PHC2208_n2195 (.Y(FE_PHN2208_n2195), 
	.A(FE_PHN3739_n2195));
   DLY4X1 FE_PHC2207_n1840 (.Y(FE_PHN2207_n1840), 
	.A(FE_PHN3722_n1840));
   DLY4X1 FE_PHC2206_n1444 (.Y(FE_PHN2206_n1444), 
	.A(FE_PHN3731_n1444));
   DLY4X1 FE_PHC2205_n1492 (.Y(FE_PHN2205_n1492), 
	.A(FE_PHN3827_n1492));
   DLY4X1 FE_PHC2204_n2129 (.Y(FE_PHN2204_n2129), 
	.A(FE_PHN3707_n2129));
   DLY4X1 FE_PHC2203_n1871 (.Y(FE_PHN2203_n1871), 
	.A(FE_PHN3758_n1871));
   DLY4X1 FE_PHC2202_n2082 (.Y(FE_PHN2202_n2082), 
	.A(FE_PHN3900_n2082));
   DLY4X1 FE_PHC2201_n2193 (.Y(FE_PHN2201_n2193), 
	.A(FE_PHN3628_n2193));
   DLY4X1 FE_PHC2200_n1440 (.Y(FE_PHN2200_n1440), 
	.A(n1440));
   DLY4X1 FE_PHC2199_n2059 (.Y(FE_PHN2199_n2059), 
	.A(FE_PHN3691_n2059));
   DLY4X1 FE_PHC2198_n1679 (.Y(FE_PHN2198_n1679), 
	.A(FE_PHN3652_n1679));
   DLY4X1 FE_PHC2197_n1729 (.Y(FE_PHN2197_n1729), 
	.A(FE_PHN3768_n1729));
   DLY4X1 FE_PHC2196_n1834 (.Y(FE_PHN2196_n1834), 
	.A(FE_PHN3654_n1834));
   DLY4X1 FE_PHC2195_n2256 (.Y(FE_PHN2195_n2256), 
	.A(FE_PHN4720_n2256));
   DLY4X1 FE_PHC2194_n2285 (.Y(FE_PHN2194_n2285), 
	.A(FE_PHN4034_n2285));
   DLY4X1 FE_PHC2193_n2261 (.Y(FE_PHN2193_n2261), 
	.A(n2261));
   DLY4X1 FE_PHC2192_n1804 (.Y(FE_PHN2192_n1804), 
	.A(FE_PHN3932_n1804));
   DLY4X1 FE_PHC2191_n1482 (.Y(FE_PHN2191_n1482), 
	.A(FE_PHN3625_n1482));
   DLY4X1 FE_PHC2190_n1420 (.Y(FE_PHN2190_n1420), 
	.A(FE_PHN4160_n1420));
   DLY4X1 FE_PHC2189_n1905 (.Y(FE_PHN2189_n1905), 
	.A(n1905));
   DLY4X1 FE_PHC2188_n2054 (.Y(FE_PHN2188_n2054), 
	.A(FE_PHN3734_n2054));
   DLY4X1 FE_PHC2187_n2120 (.Y(FE_PHN2187_n2120), 
	.A(n2120));
   DLY4X1 FE_PHC2186_n2197 (.Y(FE_PHN2186_n2197), 
	.A(n2197));
   DLY4X1 FE_PHC2185_n1820 (.Y(FE_PHN2185_n1820), 
	.A(FE_PHN4565_n1820));
   DLY4X1 FE_PHC2184_n2242 (.Y(FE_PHN2184_n2242), 
	.A(FE_PHN3740_n2242));
   DLY4X1 FE_PHC2183_n1760 (.Y(FE_PHN2183_n1760), 
	.A(FE_PHN3761_n1760));
   DLY4X1 FE_PHC2182_n2282 (.Y(FE_PHN2182_n2282), 
	.A(n2282));
   DLY4X1 FE_PHC2181_n1773 (.Y(FE_PHN2181_n1773), 
	.A(FE_PHN4123_n1773));
   DLY4X1 FE_PHC2180_n2136 (.Y(FE_PHN2180_n2136), 
	.A(FE_PHN3672_n2136));
   DLY4X1 FE_PHC2179_n1497 (.Y(FE_PHN2179_n1497), 
	.A(FE_PHN3879_n1497));
   DLY4X1 FE_PHC2178_n2212 (.Y(FE_PHN2178_n2212), 
	.A(FE_PHN3629_n2212));
   DLY4X1 FE_PHC2177_n2200 (.Y(FE_PHN2177_n2200), 
	.A(FE_PHN3682_n2200));
   DLY4X1 FE_PHC2176_n2288 (.Y(FE_PHN2176_n2288), 
	.A(FE_PHN3717_n2288));
   DLY4X1 FE_PHC2175_n1722 (.Y(FE_PHN2175_n1722), 
	.A(FE_PHN3698_n1722));
   DLY4X1 FE_PHC2174_n1847 (.Y(FE_PHN2174_n1847), 
	.A(n1847));
   DLY4X1 FE_PHC2173_n1827 (.Y(FE_PHN2173_n1827), 
	.A(FE_PHN4861_n1827));
   DLY4X1 FE_PHC2172_n1705 (.Y(FE_PHN2172_n1705), 
	.A(FE_PHN3769_n1705));
   DLY4X1 FE_PHC2171_n1864 (.Y(FE_PHN2171_n1864), 
	.A(FE_PHN3690_n1864));
   DLY4X1 FE_PHC2170_n1446 (.Y(FE_PHN2170_n1446), 
	.A(FE_PHN3666_n1446));
   DLY4X1 FE_PHC2169_n1789 (.Y(FE_PHN2169_n1789), 
	.A(FE_PHN3948_n1789));
   DLY4X1 FE_PHC2168_n2190 (.Y(FE_PHN2168_n2190), 
	.A(FE_PHN3677_n2190));
   DLY4X1 FE_PHC2167_n1669 (.Y(FE_PHN2167_n1669), 
	.A(n1669));
   DLY4X1 FE_PHC2166_n1759 (.Y(FE_PHN2166_n1759), 
	.A(FE_PHN3892_n1759));
   DLY4X1 FE_PHC2165_n1715 (.Y(FE_PHN2165_n1715), 
	.A(FE_PHN3964_n1715));
   DLY4X1 FE_PHC2164_n1406 (.Y(FE_PHN2164_n1406), 
	.A(FE_PHN3753_n1406));
   DLY4X1 FE_PHC2163_n1887 (.Y(FE_PHN2163_n1887), 
	.A(FE_PHN4721_n1887));
   DLY4X1 FE_PHC2162_n2070 (.Y(FE_PHN2162_n2070), 
	.A(FE_PHN3664_n2070));
   DLY4X1 FE_PHC2161_n2181 (.Y(FE_PHN2161_n2181), 
	.A(n2181));
   DLY4X1 FE_PHC2160_n1850 (.Y(FE_PHN2160_n1850), 
	.A(FE_PHN3981_n1850));
   DLY4X1 FE_PHC2159_n2210 (.Y(FE_PHN2159_n2210), 
	.A(FE_PHN3814_n2210));
   DLY4X1 FE_PHC2158_n1904 (.Y(FE_PHN2158_n1904), 
	.A(FE_PHN3689_n1904));
   DLY4X1 FE_PHC2157_n2099 (.Y(FE_PHN2157_n2099), 
	.A(FE_PHN3708_n2099));
   DLY4X1 FE_PHC2156_n1714 (.Y(FE_PHN2156_n1714), 
	.A(FE_PHN3857_n1714));
   DLY4X1 FE_PHC2155_n2096 (.Y(FE_PHN2155_n2096), 
	.A(FE_PHN3996_n2096));
   DLY4X1 FE_PHC2154_n1489 (.Y(FE_PHN2154_n1489), 
	.A(FE_PHN3835_n1489));
   DLY4X1 FE_PHC2153_n1724 (.Y(FE_PHN2153_n1724), 
	.A(FE_PHN3619_n1724));
   DLY4X1 FE_PHC2152_n2163 (.Y(FE_PHN2152_n2163), 
	.A(FE_PHN4166_n2163));
   DLY4X1 FE_PHC2151_n1704 (.Y(FE_PHN2151_n1704), 
	.A(FE_PHN4007_n1704));
   DLY4X1 FE_PHC2150_n1774 (.Y(FE_PHN2150_n1774), 
	.A(FE_PHN3733_n1774));
   DLY4X1 FE_PHC2149_n1835 (.Y(FE_PHN2149_n1835), 
	.A(FE_PHN3824_n1835));
   DLY4X1 FE_PHC2148_n1848 (.Y(FE_PHN2148_n1848), 
	.A(FE_PHN3634_n1848));
   DLY4X1 FE_PHC2147_n2204 (.Y(FE_PHN2147_n2204), 
	.A(FE_PHN3711_n2204));
   DLY4X1 FE_PHC2146_n2237 (.Y(FE_PHN2146_n2237), 
	.A(FE_PHN4021_n2237));
   DLY4X1 FE_PHC2145_n2142 (.Y(FE_PHN2145_n2142), 
	.A(FE_PHN3930_n2142));
   DLY4X1 FE_PHC2144_n2160 (.Y(FE_PHN2144_n2160), 
	.A(FE_PHN3729_n2160));
   DLY4X1 FE_PHC2143_n1802 (.Y(FE_PHN2143_n1802), 
	.A(FE_PHN3929_n1802));
   DLY4X1 FE_PHC2142_n1656 (.Y(FE_PHN2142_n1656), 
	.A(FE_PHN3710_n1656));
   DLY4X1 FE_PHC2141_n1397 (.Y(FE_PHN2141_n1397), 
	.A(FE_PHN3922_n1397));
   DLY4X1 FE_PHC2140_n2175 (.Y(FE_PHN2140_n2175), 
	.A(FE_PHN3701_n2175));
   DLY4X1 FE_PHC2139_n2273 (.Y(FE_PHN2139_n2273), 
	.A(n2273));
   DLY4X1 FE_PHC2138_n2121 (.Y(FE_PHN2138_n2121), 
	.A(FE_PHN3621_n2121));
   DLY4X1 FE_PHC2137_n2206 (.Y(FE_PHN2137_n2206), 
	.A(FE_PHN3680_n2206));
   DLY4X1 FE_PHC2136_n1825 (.Y(FE_PHN2136_n1825), 
	.A(FE_PHN4235_n1825));
   DLY4X1 FE_PHC2135_n1653 (.Y(FE_PHN2135_n1653), 
	.A(FE_PHN3661_n1653));
   DLY4X1 FE_PHC2134_n1846 (.Y(FE_PHN2134_n1846), 
	.A(FE_PHN3974_n1846));
   DLY4X1 FE_PHC2133_n1424 (.Y(FE_PHN2133_n1424), 
	.A(FE_PHN3713_n1424));
   DLY4X1 FE_PHC2132_n2141 (.Y(FE_PHN2132_n2141), 
	.A(FE_PHN3705_n2141));
   DLY4X1 FE_PHC2131_n1442 (.Y(FE_PHN2131_n1442), 
	.A(FE_PHN3697_n1442));
   DLY4X1 FE_PHC2130_n1849 (.Y(FE_PHN2130_n1849), 
	.A(FE_PHN3696_n1849));
   DLY4X1 FE_PHC2129_n2137 (.Y(FE_PHN2129_n2137), 
	.A(FE_PHN3617_n2137));
   DLY4X1 FE_PHC2128_n1733 (.Y(FE_PHN2128_n1733), 
	.A(FE_PHN3685_n1733));
   DLY4X1 FE_PHC2127_n2081 (.Y(FE_PHN2127_n2081), 
	.A(FE_PHN4655_n2081));
   DLY4X1 FE_PHC2126_n2196 (.Y(FE_PHN2126_n2196), 
	.A(FE_PHN3694_n2196));
   DLY4X1 FE_PHC2125_n1894 (.Y(FE_PHN2125_n1894), 
	.A(FE_PHN3822_n1894));
   DLY4X1 FE_PHC2124_n1452 (.Y(FE_PHN2124_n1452), 
	.A(FE_PHN3668_n1452));
   DLY4X1 FE_PHC2123_n2218 (.Y(FE_PHN2123_n2218), 
	.A(FE_PHN3724_n2218));
   DLY4X1 FE_PHC2122_n1718 (.Y(FE_PHN2122_n1718), 
	.A(FE_PHN3623_n1718));
   DLY4X1 FE_PHC2121_n1486 (.Y(FE_PHN2121_n1486), 
	.A(FE_PHN3795_n1486));
   DLY4X1 FE_PHC2120_n1692 (.Y(FE_PHN2120_n1692), 
	.A(FE_PHN3676_n1692));
   DLY4X1 FE_PHC2119_n2259 (.Y(FE_PHN2119_n2259), 
	.A(FE_PHN3765_n2259));
   DLY4X1 FE_PHC2118_n1878 (.Y(FE_PHN2118_n1878), 
	.A(FE_PHN3615_n1878));
   DLY4X1 FE_PHC2117_n1826 (.Y(FE_PHN2117_n1826), 
	.A(FE_PHN4524_n1826));
   DLY4X1 FE_PHC2116_n1690 (.Y(FE_PHN2116_n1690), 
	.A(n1690));
   DLY4X1 FE_PHC2115_n2132 (.Y(FE_PHN2115_n2132), 
	.A(FE_PHN3836_n2132));
   DLY4X1 FE_PHC2114_n2251 (.Y(FE_PHN2114_n2251), 
	.A(FE_PHN3728_n2251));
   DLY4X1 FE_PHC2113_n2146 (.Y(FE_PHN2113_n2146), 
	.A(FE_PHN3727_n2146));
   DLY4X1 FE_PHC2112_n1491 (.Y(FE_PHN2112_n1491), 
	.A(FE_PHN3907_n1491));
   DLY4X1 FE_PHC2111_n1818 (.Y(FE_PHN2111_n1818), 
	.A(FE_PHN3681_n1818));
   DLY4X1 FE_PHC2110_n1880 (.Y(FE_PHN2110_n1880), 
	.A(FE_PHN3815_n1880));
   DLY4X1 FE_PHC2109_n2158 (.Y(FE_PHN2109_n2158), 
	.A(FE_PHN3662_n2158));
   DLY4X1 FE_PHC2108_n2068 (.Y(FE_PHN2108_n2068), 
	.A(FE_PHN3861_n2068));
   DLY4X1 FE_PHC2107_n1450 (.Y(FE_PHN2107_n1450), 
	.A(FE_PHN3622_n1450));
   DLY4X1 FE_PHC2106_n1666 (.Y(FE_PHN2106_n1666), 
	.A(FE_PHN3645_n1666));
   DLY4X1 FE_PHC2105_n1852 (.Y(FE_PHN2105_n1852), 
	.A(FE_PHN3878_n1852));
   DLY4X1 FE_PHC2104_n1417 (.Y(FE_PHN2104_n1417), 
	.A(FE_PHN3838_n1417));
   DLY4X1 FE_PHC2103_n1487 (.Y(FE_PHN2103_n1487), 
	.A(FE_PHN3688_n1487));
   DLY4X1 FE_PHC2102_n1713 (.Y(FE_PHN2102_n1713), 
	.A(FE_PHN3643_n1713));
   DLY4X1 FE_PHC2101_n2062 (.Y(FE_PHN2101_n2062), 
	.A(FE_PHN3916_n2062));
   DLY4X1 FE_PHC2100_n1717 (.Y(FE_PHN2100_n1717), 
	.A(FE_PHN3616_n1717));
   DLY4X1 FE_PHC2099_n1855 (.Y(FE_PHN2099_n1855), 
	.A(FE_PHN3841_n1855));
   DLY4X1 FE_PHC2098_n1422 (.Y(FE_PHN2098_n1422), 
	.A(FE_PHN3687_n1422));
   DLY4X1 FE_PHC2097_n1891 (.Y(FE_PHN2097_n1891), 
	.A(FE_PHN3614_n1891));
   DLY4X1 FE_PHC2096_n1814 (.Y(FE_PHN2096_n1814), 
	.A(FE_PHN3686_n1814));
   DLY4X1 FE_PHC2095_n1426 (.Y(FE_PHN2095_n1426), 
	.A(n1426));
   DLY4X1 FE_PHC2094_n2168 (.Y(FE_PHN2094_n2168), 
	.A(FE_PHN3915_n2168));
   DLY4X1 FE_PHC2093_n2215 (.Y(FE_PHN2093_n2215), 
	.A(FE_PHN3618_n2215));
   DLY4X1 FE_PHC2092_n1833 (.Y(FE_PHN2092_n1833), 
	.A(FE_PHN3656_n1833));
   DLY4X1 FE_PHC2091_n1407 (.Y(FE_PHN2091_n1407), 
	.A(FE_PHN4182_n1407));
   DLY4X1 FE_PHC2090_n2152 (.Y(FE_PHN2090_n2152), 
	.A(FE_PHN3644_n2152));
   DLY4X1 FE_PHC2089_n1706 (.Y(FE_PHN2089_n1706), 
	.A(FE_PHN3669_n1706));
   DLY4X1 FE_PHC2088_n2284 (.Y(FE_PHN2088_n2284), 
	.A(FE_PHN3663_n2284));
   DLY4X1 FE_PHC2087_n1425 (.Y(FE_PHN2087_n1425), 
	.A(FE_PHN3651_n1425));
   DLY4X1 FE_PHC2086_n2198 (.Y(FE_PHN2086_n2198), 
	.A(FE_PHN3754_n2198));
   DLY4X1 FE_PHC2085_n1405 (.Y(FE_PHN2085_n1405), 
	.A(FE_PHN3638_n1405));
   DLY4X1 FE_PHC2084_n2079 (.Y(FE_PHN2084_n2079), 
	.A(FE_PHN3778_n2079));
   DLY4X1 FE_PHC2083_n2214 (.Y(FE_PHN2083_n2214), 
	.A(FE_PHN3807_n2214));
   DLY4X1 FE_PHC2082_n1412 (.Y(FE_PHN2082_n1412), 
	.A(FE_PHN3650_n1412));
   DLY4X1 FE_PHC2081_n1710 (.Y(FE_PHN2081_n1710), 
	.A(FE_PHN3854_n1710));
   DLY4X1 FE_PHC2080_n1499 (.Y(FE_PHN2080_n1499), 
	.A(FE_PHN3842_n1499));
   DLY4X1 FE_PHC2079_n1496 (.Y(FE_PHN2079_n1496), 
	.A(FE_PHN4265_n1496));
   DLY4X1 FE_PHC2078_n1873 (.Y(FE_PHN2078_n1873), 
	.A(FE_PHN3837_n1873));
   DLY4X1 FE_PHC2077_n1423 (.Y(FE_PHN2077_n1423), 
	.A(FE_PHN3647_n1423));
   DLY4X1 FE_PHC2076_n2105 (.Y(FE_PHN2076_n2105), 
	.A(FE_PHN3642_n2105));
   DLY4X1 FE_PHC2075_n1762 (.Y(FE_PHN2075_n1762), 
	.A(FE_PHN3867_n1762));
   DLY4X1 FE_PHC2074_n2089 (.Y(FE_PHN2074_n2089), 
	.A(FE_PHN3791_n2089));
   DLY4X1 FE_PHC2073_n1678 (.Y(FE_PHN2073_n1678), 
	.A(FE_PHN3648_n1678));
   DLY4X1 FE_PHC2072_n2286 (.Y(FE_PHN2072_n2286), 
	.A(FE_PHN3893_n2286));
   DLY4X1 FE_PHC2071_n2138 (.Y(FE_PHN2071_n2138), 
	.A(FE_PHN4458_n2138));
   DLY4X1 FE_PHC2070_n2211 (.Y(FE_PHN2070_n2211), 
	.A(FE_PHN3953_n2211));
   DLY4X1 FE_PHC2069_n1829 (.Y(FE_PHN2069_n1829), 
	.A(FE_PHN3875_n1829));
   DLY4X1 FE_PHC2068_n1753 (.Y(FE_PHN2068_n1753), 
	.A(n1753));
   DLY4X1 FE_PHC2067_n2243 (.Y(FE_PHN2067_n2243), 
	.A(FE_PHN3908_n2243));
   DLY4X1 FE_PHC2066_n1498 (.Y(FE_PHN2066_n1498), 
	.A(FE_PHN3844_n1498));
   DLY4X1 FE_PHC2065_n1796 (.Y(FE_PHN2065_n1796), 
	.A(FE_PHN3613_n1796));
   DLY4X1 FE_PHC2064_n2246 (.Y(FE_PHN2064_n2246), 
	.A(FE_PHN3936_n2246));
   DLY4X1 FE_PHC2063_n1712 (.Y(FE_PHN2063_n1712), 
	.A(FE_PHN3641_n1712));
   DLY4X1 FE_PHC2062_n1661 (.Y(FE_PHN2062_n1661), 
	.A(FE_PHN3611_n1661));
   DLY4X1 FE_PHC2061_n1691 (.Y(FE_PHN2061_n1691), 
	.A(FE_PHN3851_n1691));
   DLY4X1 FE_PHC2060_n1490 (.Y(FE_PHN2060_n1490), 
	.A(FE_PHN3834_n1490));
   DLY4X1 FE_PHC2059_n1459 (.Y(FE_PHN2059_n1459), 
	.A(FE_PHN3921_n1459));
   DLY4X1 FE_PHC2058_n2199 (.Y(FE_PHN2058_n2199), 
	.A(FE_PHN3847_n2199));
   DLY4X1 FE_PHC2057_n2088 (.Y(FE_PHN2057_n2088), 
	.A(FE_PHN3863_n2088));
   DLY4X1 FE_PHC2056_n1764 (.Y(FE_PHN2056_n1764), 
	.A(FE_PHN3665_n1764));
   DLY4X1 FE_PHC2055_n1763 (.Y(FE_PHN2055_n1763), 
	.A(FE_PHN3612_n1763));
   DLY4X1 FE_PHC2054_n1771 (.Y(FE_PHN2054_n1771), 
	.A(FE_PHN3631_n1771));
   DLY4X1 FE_PHC2053_n2044 (.Y(FE_PHN2053_n2044), 
	.A(FE_PHN3763_n2044));
   DLY4X1 FE_PHC2052_n2221 (.Y(FE_PHN2052_n2221), 
	.A(FE_PHN4060_n2221));
   DLY4X1 FE_PHC2051_n1805 (.Y(FE_PHN2051_n1805), 
	.A(FE_PHN3787_n1805));
   DLY4X1 FE_PHC2050_n1687 (.Y(FE_PHN2050_n1687), 
	.A(FE_PHN3671_n1687));
   DLY4X1 FE_PHC2049_n1885 (.Y(FE_PHN2049_n1885), 
	.A(FE_PHN4190_n1885));
   DLY4X1 FE_PHC2048_n2235 (.Y(FE_PHN2048_n2235), 
	.A(FE_PHN3626_n2235));
   DLY4X1 FE_PHC2047_n2104 (.Y(FE_PHN2047_n2104), 
	.A(n2104));
   DLY4X1 FE_PHC2046_n1416 (.Y(FE_PHN2046_n1416), 
	.A(FE_PHN3633_n1416));
   DLY4X1 FE_PHC2045_n2073 (.Y(FE_PHN2045_n2073), 
	.A(FE_PHN3640_n2073));
   DLY4X1 FE_PHC2044_n1732 (.Y(FE_PHN2044_n1732), 
	.A(n1732));
   DLY4X1 FE_PHC2043_n1769 (.Y(FE_PHN2043_n1769), 
	.A(FE_PHN3755_n1769));
   DLY4X1 FE_PHC2042_n2069 (.Y(FE_PHN2042_n2069), 
	.A(FE_PHN3743_n2069));
   DLY4X1 FE_PHC2041_n2098 (.Y(FE_PHN2041_n2098), 
	.A(FE_PHN3737_n2098));
   DLY4X1 FE_PHC2040_n2092 (.Y(FE_PHN2040_n2092), 
	.A(FE_PHN3674_n2092));
   DLY4X1 FE_PHC2039_n1511 (.Y(FE_PHN2039_n1511), 
	.A(FE_PHN3735_n1511));
   DLY4X1 FE_PHC2038_n2393 (.Y(FE_PHN2038_n2393), 
	.A(FE_PHN5053_n2393));
   DLY4X1 FE_PHC2036_n2394 (.Y(FE_PHN2036_n2394), 
	.A(FE_PHN5042_n2394));
   DLY4X1 FE_PHC2009_n1799 (.Y(FE_PHN2009_n1799), 
	.A(FE_PHN4143_n1799));
   DLY4X1 FE_PHC2008_n1786 (.Y(FE_PHN2008_n1786), 
	.A(FE_PHN3865_n1786));
   DLY4X1 FE_PHC2007_keymem_sboxw_13_ (.Y(sboxw[13]), 
	.A(FE_PHN2007_keymem_sboxw_13_));
   DLY4X1 FE_PHC2006_keymem_sboxw_5_ (.Y(FE_PHN2006_keymem_sboxw_5_), 
	.A(sboxw[5]));
   DLY4X1 FE_PHC2005_keymem_sboxw_20_ (.Y(FE_PHN2005_keymem_sboxw_20_), 
	.A(sboxw[20]));
   DLY4X1 FE_PHC2004_keymem_sboxw_12_ (.Y(FE_PHN2004_keymem_sboxw_12_), 
	.A(sboxw[12]));
   DLY4X1 FE_PHC2003_keymem_sboxw_4_ (.Y(FE_PHN2003_keymem_sboxw_4_), 
	.A(sboxw[4]));
   DLY4X1 FE_PHC2002_keymem_sboxw_11_ (.Y(sboxw[11]), 
	.A(FE_PHN2002_keymem_sboxw_11_));
   DLY4X1 FE_PHC2001_keymem_sboxw_8_ (.Y(FE_PHN2001_keymem_sboxw_8_), 
	.A(sboxw[8]));
   DLY4X1 FE_PHC2000_keymem_sboxw_3_ (.Y(sboxw[3]), 
	.A(FE_PHN2000_keymem_sboxw_3_));
   DLY4X1 FE_PHC1998_keymem_sboxw_17_ (.Y(FE_PHN1998_keymem_sboxw_17_), 
	.A(sboxw[17]));
   DLY4X1 FE_PHC1997_keymem_sboxw_16_ (.Y(sboxw[16]), 
	.A(FE_PHN1997_keymem_sboxw_16_));
   DLY4X1 FE_PHC1992_keymem_sboxw_19_ (.Y(sboxw[19]), 
	.A(FE_PHN1992_keymem_sboxw_19_));
   DLY4X1 FE_PHC1991_keymem_sboxw_9_ (.Y(sboxw[9]), 
	.A(FE_PHN1991_keymem_sboxw_9_));
   DLY4X1 FE_PHC1989_rcon_reg_6_ (.Y(FE_PHN1989_rcon_reg_6_), 
	.A(rcon_reg[6]));
   DLY4X1 FE_PHC1974_keymem_sboxw_14_ (.Y(sboxw[14]), 
	.A(FE_PHN1974_keymem_sboxw_14_));
   DLY4X1 FE_PHC1972_keymem_sboxw_15_ (.Y(sboxw[15]), 
	.A(FE_PHN1972_keymem_sboxw_15_));
   DLY4X1 FE_PHC1969_keymem_sboxw_23_ (.Y(sboxw[23]), 
	.A(FE_PHN1969_keymem_sboxw_23_));
   DLY4X1 FE_PHC1965_keymem_sboxw_22_ (.Y(FE_PHN1965_keymem_sboxw_22_), 
	.A(sboxw[22]));
   DLY4X1 FE_PHC1962_keymem_sboxw_10_ (.Y(FE_PHN1962_keymem_sboxw_10_), 
	.A(sboxw[10]));
   DLY4X1 FE_PHC1959_keymem_sboxw_0_ (.Y(FE_PHN1959_keymem_sboxw_0_), 
	.A(sboxw[0]));
   DLY4X1 FE_PHC1958_keymem_sboxw_18_ (.Y(FE_PHN1958_keymem_sboxw_18_), 
	.A(sboxw[18]));
   DLY4X1 FE_PHC1957_keymem_sboxw_1_ (.Y(sboxw[1]), 
	.A(FE_PHN1957_keymem_sboxw_1_));
   DLY4X1 FE_PHC1930_key_mem_1082_ (.Y(FE_PHN1930_key_mem_1082_), 
	.A(key_mem[1082]));
   DLY4X1 FE_PHC1917_key_mem_1207_ (.Y(FE_PHN1917_key_mem_1207_), 
	.A(key_mem[1207]));
   DLY4X1 FE_PHC1905_key_mem_1046_ (.Y(FE_PHN1905_key_mem_1046_), 
	.A(key_mem[1046]));
   DLY4X1 FE_PHC1899_key_mem_1272_ (.Y(FE_PHN1899_key_mem_1272_), 
	.A(key_mem[1272]));
   DLY4X1 FE_PHC1894_key_mem_1044_ (.Y(FE_PHN1894_key_mem_1044_), 
	.A(key_mem[1044]));
   DLY4X1 FE_PHC1893_key_mem_1101_ (.Y(FE_PHN1893_key_mem_1101_), 
	.A(key_mem[1101]));
   DLY4X1 FE_PHC1892_key_mem_1029_ (.Y(FE_PHN1892_key_mem_1029_), 
	.A(key_mem[1029]));
   DLY4X1 FE_PHC1891_key_mem_1068_ (.Y(FE_PHN1891_key_mem_1068_), 
	.A(key_mem[1068]));
   DLY4X1 FE_PHC1889_key_mem_1071_ (.Y(FE_PHN1889_key_mem_1071_), 
	.A(key_mem[1071]));
   DLY4X1 FE_PHC1888_key_mem_1039_ (.Y(FE_PHN1888_key_mem_1039_), 
	.A(key_mem[1039]));
   DLY4X1 FE_PHC1887_key_mem_1100_ (.Y(FE_PHN1887_key_mem_1100_), 
	.A(key_mem[1100]));
   DLY4X1 FE_PHC1885_key_mem_1114_ (.Y(FE_PHN1885_key_mem_1114_), 
	.A(key_mem[1114]));
   DLY4X1 FE_PHC1884_key_mem_1151_ (.Y(FE_PHN1884_key_mem_1151_), 
	.A(key_mem[1151]));
   DLY4X1 FE_PHC1883_key_mem_1153_ (.Y(FE_PHN1883_key_mem_1153_), 
	.A(key_mem[1153]));
   DLY4X1 FE_PHC1882_key_mem_1025_ (.Y(FE_PHN1882_key_mem_1025_), 
	.A(key_mem[1025]));
   DLY4X1 FE_PHC1881_key_mem_1040_ (.Y(FE_PHN1881_key_mem_1040_), 
	.A(key_mem[1040]));
   DLY4X1 FE_PHC1880_key_mem_1045_ (.Y(FE_PHN1880_key_mem_1045_), 
	.A(key_mem[1045]));
   DLY4X1 FE_PHC1879_key_mem_688_ (.Y(FE_PHN1879_key_mem_688_), 
	.A(key_mem[688]));
   DLY4X1 FE_PHC1878_n1167 (.Y(FE_PHN1878_n1167), 
	.A(FE_PHN4723_n1167));
   DLY4X1 FE_PHC1877_key_mem_1255_ (.Y(FE_PHN1877_key_mem_1255_), 
	.A(key_mem[1255]));
   DLY4X1 FE_PHC1876_key_mem_1049_ (.Y(FE_PHN1876_key_mem_1049_), 
	.A(key_mem[1049]));
   DLY4X1 FE_PHC1874_key_mem_1143_ (.Y(FE_PHN1874_key_mem_1143_), 
	.A(key_mem[1143]));
   DLY4X1 FE_PHC1873_key_mem_1061_ (.Y(FE_PHN1873_key_mem_1061_), 
	.A(key_mem[1061]));
   DLY4X1 FE_PHC1872_key_mem_1060_ (.Y(FE_PHN1872_key_mem_1060_), 
	.A(key_mem[1060]));
   DLY4X1 FE_PHC1871_key_mem_1106_ (.Y(FE_PHN1871_key_mem_1106_), 
	.A(key_mem[1106]));
   DLY4X1 FE_PHC1870_key_mem_1138_ (.Y(FE_PHN1870_key_mem_1138_), 
	.A(key_mem[1138]));
   DLY4X1 FE_PHC1869_key_mem_1088_ (.Y(FE_PHN1869_key_mem_1088_), 
	.A(key_mem[1088]));
   DLY4X1 FE_PHC1868_key_mem_1053_ (.Y(FE_PHN1868_key_mem_1053_), 
	.A(key_mem[1053]));
   DLY4X1 FE_PHC1867_key_mem_1069_ (.Y(FE_PHN1867_key_mem_1069_), 
	.A(key_mem[1069]));
   DLY4X1 FE_PHC1866_key_mem_1078_ (.Y(FE_PHN1866_key_mem_1078_), 
	.A(key_mem[1078]));
   DLY4X1 FE_PHC1864_key_mem_1055_ (.Y(FE_PHN1864_key_mem_1055_), 
	.A(key_mem[1055]));
   DLY4X1 FE_PHC1863_key_mem_1094_ (.Y(FE_PHN1863_key_mem_1094_), 
	.A(key_mem[1094]));
   DLY4X1 FE_PHC1862_key_mem_1030_ (.Y(FE_PHN1862_key_mem_1030_), 
	.A(key_mem[1030]));
   DLY4X1 FE_PHC1861_key_mem_1072_ (.Y(FE_PHN1861_key_mem_1072_), 
	.A(key_mem[1072]));
   DLY4X1 FE_PHC1860_key_mem_1112_ (.Y(FE_PHN1860_key_mem_1112_), 
	.A(key_mem[1112]));
   DLY4X1 FE_PHC1859_key_mem_1099_ (.Y(FE_PHN1859_key_mem_1099_), 
	.A(key_mem[1099]));
   DLY4X1 FE_PHC1858_key_mem_1144_ (.Y(FE_PHN1858_key_mem_1144_), 
	.A(key_mem[1144]));
   DLY4X1 FE_PHC1857_key_mem_1083_ (.Y(FE_PHN1857_key_mem_1083_), 
	.A(key_mem[1083]));
   DLY4X1 FE_PHC1856_key_mem_1085_ (.Y(FE_PHN1856_key_mem_1085_), 
	.A(key_mem[1085]));
   DLY4X1 FE_PHC1855_key_mem_1103_ (.Y(FE_PHN1855_key_mem_1103_), 
	.A(key_mem[1103]));
   DLY4X1 FE_PHC1854_key_mem_1127_ (.Y(FE_PHN1854_key_mem_1127_), 
	.A(key_mem[1127]));
   DLY4X1 FE_PHC1853_key_mem_1028_ (.Y(FE_PHN1853_key_mem_1028_), 
	.A(key_mem[1028]));
   DLY4X1 FE_PHC1852_key_mem_1064_ (.Y(FE_PHN1852_key_mem_1064_), 
	.A(key_mem[1064]));
   DLY4X1 FE_PHC1851_key_mem_349_ (.Y(FE_PHN1851_key_mem_349_), 
	.A(key_mem[349]));
   DLY4X1 FE_PHC1850_key_mem_1121_ (.Y(FE_PHN1850_key_mem_1121_), 
	.A(key_mem[1121]));
   DLY4X1 FE_PHC1849_key_mem_376_ (.Y(FE_PHN1849_key_mem_376_), 
	.A(key_mem[376]));
   DLY4X1 FE_PHC1848_key_mem_647_ (.Y(FE_PHN1848_key_mem_647_), 
	.A(key_mem[647]));
   DLY4X1 FE_PHC1847_n1162 (.Y(FE_PHN1847_n1162), 
	.A(n1162));
   DLY4X1 FE_PHC1846_key_mem_1142_ (.Y(FE_PHN1846_key_mem_1142_), 
	.A(key_mem[1142]));
   DLY4X1 FE_PHC1844_key_mem_352_ (.Y(FE_PHN1844_key_mem_352_), 
	.A(key_mem[352]));
   DLY4X1 FE_PHC1843_key_mem_1116_ (.Y(FE_PHN1843_key_mem_1116_), 
	.A(key_mem[1116]));
   DLY4X1 FE_PHC1841_key_mem_1092_ (.Y(FE_PHN1841_key_mem_1092_), 
	.A(key_mem[1092]));
   DLY4X1 FE_PHC1840_key_mem_1041_ (.Y(FE_PHN1840_key_mem_1041_), 
	.A(key_mem[1041]));
   DLY4X1 FE_PHC1839_key_mem_1059_ (.Y(FE_PHN1839_key_mem_1059_), 
	.A(key_mem[1059]));
   DLY4X1 FE_PHC1837_n2267 (.Y(FE_PHN1837_n2267), 
	.A(FE_PHN4393_n2267));
   DLY4X1 FE_PHC1835_key_mem_1084_ (.Y(FE_PHN1835_key_mem_1084_), 
	.A(key_mem[1084]));
   DLY4X1 FE_PHC1834_key_mem_1311_ (.Y(FE_PHN1834_key_mem_1311_), 
	.A(key_mem[1311]));
   DLY4X1 FE_PHC1833_key_mem_1043_ (.Y(FE_PHN1833_key_mem_1043_), 
	.A(key_mem[1043]));
   DLY4X1 FE_PHC1832_key_mem_1057_ (.Y(FE_PHN1832_key_mem_1057_), 
	.A(key_mem[1057]));
   DLY4X1 FE_PHC1831_key_mem_724_ (.Y(FE_PHN1831_key_mem_724_), 
	.A(key_mem[724]));
   DLY4X1 FE_PHC1830_key_mem_1090_ (.Y(FE_PHN1830_key_mem_1090_), 
	.A(key_mem[1090]));
   DLY4X1 FE_PHC1829_key_mem_1079_ (.Y(FE_PHN1829_key_mem_1079_), 
	.A(key_mem[1079]));
   DLY4X1 FE_PHC1828_key_mem_755_ (.Y(FE_PHN1828_key_mem_755_), 
	.A(key_mem[755]));
   DLY4X1 FE_PHC1827_n1181 (.Y(FE_PHN1827_n1181), 
	.A(FE_PHN4557_n1181));
   DLY4X1 FE_PHC1826_key_mem_334_ (.Y(FE_PHN1826_key_mem_334_), 
	.A(key_mem[334]));
   DLY4X1 FE_PHC1824_key_mem_738_ (.Y(FE_PHN1824_key_mem_738_), 
	.A(key_mem[738]));
   DLY4X1 FE_PHC1823_key_mem_1115_ (.Y(FE_PHN1823_key_mem_1115_), 
	.A(key_mem[1115]));
   DLY4X1 FE_PHC1822_key_mem_1133_ (.Y(FE_PHN1822_key_mem_1133_), 
	.A(key_mem[1133]));
   DLY4X1 FE_PHC1821_key_mem_1104_ (.Y(FE_PHN1821_key_mem_1104_), 
	.A(key_mem[1104]));
   DLY4X1 FE_PHC1820_key_mem_713_ (.Y(FE_PHN1820_key_mem_713_), 
	.A(key_mem[713]));
   DLY4X1 FE_PHC1819_key_mem_1140_ (.Y(FE_PHN1819_key_mem_1140_), 
	.A(key_mem[1140]));
   DLY4X1 FE_PHC1818_key_mem_1113_ (.Y(FE_PHN1818_key_mem_1113_), 
	.A(key_mem[1113]));
   DLY4X1 FE_PHC1817_key_mem_1119_ (.Y(FE_PHN1817_key_mem_1119_), 
	.A(key_mem[1119]));
   DLY4X1 FE_PHC1816_key_mem_1128_ (.Y(FE_PHN1816_key_mem_1128_), 
	.A(key_mem[1128]));
   DLY4X1 FE_PHC1814_key_mem_1150_ (.Y(FE_PHN1814_key_mem_1150_), 
	.A(key_mem[1150]));
   DLY4X1 FE_PHC1813_key_mem_1066_ (.Y(FE_PHN1813_key_mem_1066_), 
	.A(key_mem[1066]));
   DLY4X1 FE_PHC1812_n1595 (.Y(FE_PHN1812_n1595), 
	.A(n1595));
   DLY4X1 FE_PHC1811_key_mem_1036_ (.Y(FE_PHN1811_key_mem_1036_), 
	.A(key_mem[1036]));
   DLY4X1 FE_PHC1810_key_mem_1136_ (.Y(FE_PHN1810_key_mem_1136_), 
	.A(key_mem[1136]));
   DLY4X1 FE_PHC1809_key_mem_644_ (.Y(FE_PHN1809_key_mem_644_), 
	.A(key_mem[644]));
   DLY4X1 FE_PHC1808_key_mem_1148_ (.Y(FE_PHN1808_key_mem_1148_), 
	.A(key_mem[1148]));
   DLY4X1 FE_PHC1807_key_mem_360_ (.Y(FE_PHN1807_key_mem_360_), 
	.A(key_mem[360]));
   DLY4X1 FE_PHC1806_key_mem_318_ (.Y(FE_PHN1806_key_mem_318_), 
	.A(key_mem[318]));
   DLY4X1 FE_PHC1805_key_mem_1147_ (.Y(FE_PHN1805_key_mem_1147_), 
	.A(key_mem[1147]));
   DLY4X1 FE_PHC1804_key_mem_737_ (.Y(FE_PHN1804_key_mem_737_), 
	.A(key_mem[737]));
   DLY4X1 FE_PHC1803_key_mem_1118_ (.Y(FE_PHN1803_key_mem_1118_), 
	.A(key_mem[1118]));
   DLY4X1 FE_PHC1802_key_mem_285_ (.Y(FE_PHN1802_key_mem_285_), 
	.A(key_mem[285]));
   DLY4X1 FE_PHC1801_n1240 (.Y(FE_PHN1801_n1240), 
	.A(FE_PHN4369_n1240));
   DLY4X1 FE_PHC1800_key_mem_1191_ (.Y(FE_PHN1800_key_mem_1191_), 
	.A(key_mem[1191]));
   DLY4X1 FE_PHC1799_key_mem_1097_ (.Y(FE_PHN1799_key_mem_1097_), 
	.A(key_mem[1097]));
   DLY4X1 FE_PHC1798_key_mem_1076_ (.Y(FE_PHN1798_key_mem_1076_), 
	.A(key_mem[1076]));
   DLY4X1 FE_PHC1797_key_mem_661_ (.Y(FE_PHN1797_key_mem_661_), 
	.A(key_mem[661]));
   DLY4X1 FE_PHC1796_n1579 (.Y(FE_PHN1796_n1579), 
	.A(FE_PHN4551_n1579));
   DLY4X1 FE_PHC1795_key_mem_311_ (.Y(FE_PHN1795_key_mem_311_), 
	.A(key_mem[311]));
   DLY4X1 FE_PHC1794_key_mem_709_ (.Y(FE_PHN1794_key_mem_709_), 
	.A(key_mem[709]));
   DLY4X1 FE_PHC1793_key_mem_353_ (.Y(FE_PHN1793_key_mem_353_), 
	.A(key_mem[353]));
   DLY4X1 FE_PHC1792_key_mem_1169_ (.Y(FE_PHN1792_key_mem_1169_), 
	.A(key_mem[1169]));
   DLY4X1 FE_PHC1791_key_mem_1135_ (.Y(FE_PHN1791_key_mem_1135_), 
	.A(key_mem[1135]));
   DLY4X1 FE_PHC1790_key_mem_1093_ (.Y(FE_PHN1790_key_mem_1093_), 
	.A(key_mem[1093]));
   DLY4X1 FE_PHC1789_key_mem_1077_ (.Y(FE_PHN1789_key_mem_1077_), 
	.A(key_mem[1077]));
   DLY4X1 FE_PHC1788_key_mem_1037_ (.Y(FE_PHN1788_key_mem_1037_), 
	.A(key_mem[1037]));
   DLY4X1 FE_PHC1787_key_mem_1109_ (.Y(FE_PHN1787_key_mem_1109_), 
	.A(key_mem[1109]));
   DLY4X1 FE_PHC1786_key_mem_1134_ (.Y(FE_PHN1786_key_mem_1134_), 
	.A(key_mem[1134]));
   DLY4X1 FE_PHC1785_key_mem_302_ (.Y(FE_PHN1785_key_mem_302_), 
	.A(key_mem[302]));
   DLY4X1 FE_PHC1784_key_mem_1051_ (.Y(FE_PHN1784_key_mem_1051_), 
	.A(key_mem[1051]));
   DLY4X1 FE_PHC1783_key_mem_1081_ (.Y(FE_PHN1783_key_mem_1081_), 
	.A(key_mem[1081]));
   DLY4X1 FE_PHC1782_n2179 (.Y(FE_PHN1782_n2179), 
	.A(FE_PHN4260_n2179));
   DLY4X1 FE_PHC1781_key_mem_1123_ (.Y(FE_PHN1781_key_mem_1123_), 
	.A(key_mem[1123]));
   DLY4X1 FE_PHC1780_key_mem_1267_ (.Y(FE_PHN1780_key_mem_1267_), 
	.A(key_mem[1267]));
   DLY4X1 FE_PHC1779_key_mem_694_ (.Y(FE_PHN1779_key_mem_694_), 
	.A(key_mem[694]));
   DLY4X1 FE_PHC1778_key_mem_1095_ (.Y(FE_PHN1778_key_mem_1095_), 
	.A(key_mem[1095]));
   DLY4X1 FE_PHC1777_key_mem_1132_ (.Y(FE_PHN1777_key_mem_1132_), 
	.A(key_mem[1132]));
   DLY4X1 FE_PHC1776_key_mem_684_ (.Y(FE_PHN1776_key_mem_684_), 
	.A(key_mem[684]));
   DLY4X1 FE_PHC1775_key_mem_344_ (.Y(FE_PHN1775_key_mem_344_), 
	.A(key_mem[344]));
   DLY4X1 FE_PHC1774_n1266 (.Y(FE_PHN1774_n1266), 
	.A(n1266));
   DLY4X1 FE_PHC1773_key_mem_1074_ (.Y(FE_PHN1773_key_mem_1074_), 
	.A(key_mem[1074]));
   DLY4X1 FE_PHC1772_key_mem_1050_ (.Y(FE_PHN1772_key_mem_1050_), 
	.A(key_mem[1050]));
   DLY4X1 FE_PHC1771_key_mem_696_ (.Y(FE_PHN1771_key_mem_696_), 
	.A(key_mem[696]));
   DLY4X1 FE_PHC1770_key_mem_723_ (.Y(FE_PHN1770_key_mem_723_), 
	.A(key_mem[723]));
   DLY4X1 FE_PHC1769_key_mem_1054_ (.Y(FE_PHN1769_key_mem_1054_), 
	.A(key_mem[1054]));
   DLY4X1 FE_PHC1768_n2047 (.Y(FE_PHN1768_n2047), 
	.A(FE_PHN4206_n2047));
   DLY4X1 FE_PHC1767_n1257 (.Y(FE_PHN1767_n1257), 
	.A(FE_PHN4217_n1257));
   DLY4X1 FE_PHC1766_key_mem_1278_ (.Y(FE_PHN1766_key_mem_1278_), 
	.A(key_mem[1278]));
   DLY4X1 FE_PHC1765_key_mem_764_ (.Y(FE_PHN1765_key_mem_764_), 
	.A(key_mem[764]));
   DLY4X1 FE_PHC1764_key_mem_1137_ (.Y(FE_PHN1764_key_mem_1137_), 
	.A(key_mem[1137]));
   DLY4X1 FE_PHC1763_key_mem_689_ (.Y(FE_PHN1763_key_mem_689_), 
	.A(key_mem[689]));
   DLY4X1 FE_PHC1762_key_mem_1145_ (.Y(FE_PHN1762_key_mem_1145_), 
	.A(key_mem[1145]));
   DLY4X1 FE_PHC1761_key_mem_1047_ (.Y(FE_PHN1761_key_mem_1047_), 
	.A(key_mem[1047]));
   DLY4X1 FE_PHC1760_key_mem_1031_ (.Y(FE_PHN1760_key_mem_1031_), 
	.A(key_mem[1031]));
   DLY4X1 FE_PHC1759_n1668 (.Y(FE_PHN1759_n1668), 
	.A(FE_PHN4197_n1668));
   DLY4X1 FE_PHC1758_key_mem_1070_ (.Y(FE_PHN1758_key_mem_1070_), 
	.A(key_mem[1070]));
   DLY4X1 FE_PHC1757_key_mem_359_ (.Y(FE_PHN1757_key_mem_359_), 
	.A(key_mem[359]));
   DLY4X1 FE_PHC1756_key_mem_1098_ (.Y(FE_PHN1756_key_mem_1098_), 
	.A(key_mem[1098]));
   DLY4X1 FE_PHC1755_key_mem_708_ (.Y(FE_PHN1755_key_mem_708_), 
	.A(key_mem[708]));
   DLY4X1 FE_PHC1754_key_mem_351_ (.Y(FE_PHN1754_key_mem_351_), 
	.A(key_mem[351]));
   DLY4X1 FE_PHC1752_n1168 (.Y(FE_PHN1752_n1168), 
	.A(FE_PHN4432_n1168));
   DLY4X1 FE_PHC1751_key_mem_758_ (.Y(FE_PHN1751_key_mem_758_), 
	.A(key_mem[758]));
   DLY4X1 FE_PHC1750_key_mem_707_ (.Y(FE_PHN1750_key_mem_707_), 
	.A(key_mem[707]));
   DLY4X1 FE_PHC1749_key_mem_675_ (.Y(FE_PHN1749_key_mem_675_), 
	.A(key_mem[675]));
   DLY4X1 FE_PHC1748_key_mem_1141_ (.Y(FE_PHN1748_key_mem_1141_), 
	.A(key_mem[1141]));
   DLY4X1 FE_PHC1747_key_mem_682_ (.Y(FE_PHN1747_key_mem_682_), 
	.A(key_mem[682]));
   DLY4X1 FE_PHC1746_key_mem_732_ (.Y(FE_PHN1746_key_mem_732_), 
	.A(key_mem[732]));
   DLY4X1 FE_PHC1745_key_mem_1105_ (.Y(FE_PHN1745_key_mem_1105_), 
	.A(key_mem[1105]));
   DLY4X1 FE_PHC1744_key_mem_659_ (.Y(FE_PHN1744_key_mem_659_), 
	.A(key_mem[659]));
   DLY4X1 FE_PHC1743_key_mem_1058_ (.Y(FE_PHN1743_key_mem_1058_), 
	.A(key_mem[1058]));
   DLY4X1 FE_PHC1742_key_mem_328_ (.Y(FE_PHN1742_key_mem_328_), 
	.A(key_mem[328]));
   DLY4X1 FE_PHC1740_key_mem_1120_ (.Y(FE_PHN1740_key_mem_1120_), 
	.A(key_mem[1120]));
   DLY4X1 FE_PHC1739_key_mem_345_ (.Y(FE_PHN1739_key_mem_345_), 
	.A(key_mem[345]));
   DLY4X1 FE_PHC1738_key_mem_260_ (.Y(FE_PHN1738_key_mem_260_), 
	.A(key_mem[260]));
   DLY4X1 FE_PHC1737_n1895 (.Y(FE_PHN1737_n1895), 
	.A(n1895));
   DLY4X1 FE_PHC1736_n1596 (.Y(FE_PHN1736_n1596), 
	.A(n1596));
   DLY4X1 FE_PHC1735_key_mem_291_ (.Y(FE_PHN1735_key_mem_291_), 
	.A(key_mem[291]));
   DLY4X1 FE_PHC1734_key_mem_1152_ (.Y(FE_PHN1734_key_mem_1152_), 
	.A(key_mem[1152]));
   DLY4X1 FE_PHC1733_n1547 (.Y(FE_PHN1733_n1547), 
	.A(FE_PHN4020_n1547));
   DLY4X1 FE_PHC1732_n1751 (.Y(FE_PHN1732_n1751), 
	.A(FE_PHN4201_n1751));
   DLY4X1 FE_PHC1731_key_mem_693_ (.Y(FE_PHN1731_key_mem_693_), 
	.A(key_mem[693]));
   DLY4X1 FE_PHC1730_key_mem_1080_ (.Y(FE_PHN1730_key_mem_1080_), 
	.A(key_mem[1080]));
   DLY4X1 FE_PHC1729_key_mem_297_ (.Y(FE_PHN1729_key_mem_297_), 
	.A(key_mem[297]));
   DLY4X1 FE_PHC1728_n2185 (.Y(FE_PHN1728_n2185), 
	.A(FE_PHN4567_n2185));
   DLY4X1 FE_PHC1727_key_mem_269_ (.Y(FE_PHN1727_key_mem_269_), 
	.A(key_mem[269]));
   DLY4X1 FE_PHC1726_key_mem_374_ (.Y(FE_PHN1726_key_mem_374_), 
	.A(key_mem[374]));
   DLY4X1 FE_PHC1725_key_mem_348_ (.Y(FE_PHN1725_key_mem_348_), 
	.A(key_mem[348]));
   DLY4X1 FE_PHC1724_key_mem_660_ (.Y(FE_PHN1724_key_mem_660_), 
	.A(key_mem[660]));
   DLY4X1 FE_PHC1723_key_mem_759_ (.Y(FE_PHN1723_key_mem_759_), 
	.A(key_mem[759]));
   DLY4X1 FE_PHC1722_key_mem_648_ (.Y(FE_PHN1722_key_mem_648_), 
	.A(key_mem[648]));
   DLY4X1 FE_PHC1721_key_mem_704_ (.Y(FE_PHN1721_key_mem_704_), 
	.A(key_mem[704]));
   DLY4X1 FE_PHC1720_key_mem_1188_ (.Y(FE_PHN1720_key_mem_1188_), 
	.A(key_mem[1188]));
   DLY4X1 FE_PHC1719_key_mem_1042_ (.Y(FE_PHN1719_key_mem_1042_), 
	.A(key_mem[1042]));
   DLY4X1 FE_PHC1718_key_mem_721_ (.Y(FE_PHN1718_key_mem_721_), 
	.A(key_mem[721]));
   DLY4X1 FE_PHC1717_key_mem_309_ (.Y(FE_PHN1717_key_mem_309_), 
	.A(key_mem[309]));
   DLY4X1 FE_PHC1716_key_mem_324_ (.Y(FE_PHN1716_key_mem_324_), 
	.A(key_mem[324]));
   DLY4X1 FE_PHC1715_key_mem_279_ (.Y(FE_PHN1715_key_mem_279_), 
	.A(key_mem[279]));
   DLY4X1 FE_PHC1714_key_mem_341_ (.Y(FE_PHN1714_key_mem_341_), 
	.A(key_mem[341]));
   DLY4X1 FE_PHC1713_key_mem_1032_ (.Y(FE_PHN1713_key_mem_1032_), 
	.A(key_mem[1032]));
   DLY4X1 FE_PHC1712_key_mem_1075_ (.Y(FE_PHN1712_key_mem_1075_), 
	.A(key_mem[1075]));
   DLY4X1 FE_PHC1711_key_mem_256_ (.Y(FE_PHN1711_key_mem_256_), 
	.A(key_mem[256]));
   DLY4X1 FE_PHC1710_key_mem_316_ (.Y(FE_PHN1710_key_mem_316_), 
	.A(key_mem[316]));
   DLY4X1 FE_PHC1709_n1258 (.Y(FE_PHN1709_n1258), 
	.A(n1258));
   DLY4X1 FE_PHC1708_n1734 (.Y(FE_PHN1708_n1734), 
	.A(FE_PHN4419_n1734));
   DLY4X1 FE_PHC1707_key_mem_343_ (.Y(FE_PHN1707_key_mem_343_), 
	.A(key_mem[343]));
   DLY4X1 FE_PHC1706_key_mem_671_ (.Y(FE_PHN1706_key_mem_671_), 
	.A(key_mem[671]));
   DLY4X1 FE_PHC1705_n2143 (.Y(FE_PHN1705_n2143), 
	.A(FE_PHN3903_n2143));
   DLY4X1 FE_PHC1703_key_mem_258_ (.Y(FE_PHN1703_key_mem_258_), 
	.A(key_mem[258]));
   DLY4X1 FE_PHC1702_key_mem_710_ (.Y(FE_PHN1702_key_mem_710_), 
	.A(key_mem[710]));
   DLY4X1 FE_PHC1701_key_mem_1089_ (.Y(FE_PHN1701_key_mem_1089_), 
	.A(key_mem[1089]));
   DLY4X1 FE_PHC1700_key_mem_1215_ (.Y(FE_PHN1700_key_mem_1215_), 
	.A(key_mem[1215]));
   DLY4X1 FE_PHC1699_key_mem_262_ (.Y(FE_PHN1699_key_mem_262_), 
	.A(key_mem[262]));
   DLY4X1 FE_PHC1698_key_mem_698_ (.Y(FE_PHN1698_key_mem_698_), 
	.A(key_mem[698]));
   DLY4X1 FE_PHC1697_key_mem_266_ (.Y(FE_PHN1697_key_mem_266_), 
	.A(key_mem[266]));
   DLY4X1 FE_PHC1696_key_mem_680_ (.Y(FE_PHN1696_key_mem_680_), 
	.A(key_mem[680]));
   DLY4X1 FE_PHC1695_key_mem_716_ (.Y(FE_PHN1695_key_mem_716_), 
	.A(key_mem[716]));
   DLY4X1 FE_PHC1694_key_mem_673_ (.Y(FE_PHN1694_key_mem_673_), 
	.A(key_mem[673]));
   DLY4X1 FE_PHC1693_n1578 (.Y(FE_PHN1693_n1578), 
	.A(FE_PHN4045_n1578));
   DLY4X1 FE_PHC1692_key_mem_739_ (.Y(FE_PHN1692_key_mem_739_), 
	.A(key_mem[739]));
   DLY4X1 FE_PHC1691_key_mem_308_ (.Y(FE_PHN1691_key_mem_308_), 
	.A(key_mem[308]));
   DLY4X1 FE_PHC1690_key_mem_346_ (.Y(FE_PHN1690_key_mem_346_), 
	.A(key_mem[346]));
   DLY4X1 FE_PHC1689_key_mem_325_ (.Y(FE_PHN1689_key_mem_325_), 
	.A(key_mem[325]));
   DLY4X1 FE_PHC1688_key_mem_265_ (.Y(FE_PHN1688_key_mem_265_), 
	.A(key_mem[265]));
   DLY4X1 FE_PHC1687_key_mem_662_ (.Y(FE_PHN1687_key_mem_662_), 
	.A(key_mem[662]));
   DLY4X1 FE_PHC1686_n1438 (.Y(FE_PHN1686_n1438), 
	.A(FE_PHN3792_n1438));
   DLY4X1 FE_PHC1685_n1896 (.Y(FE_PHN1685_n1896), 
	.A(FE_PHN3999_n1896));
   DLY4X1 FE_PHC1684_key_mem_288_ (.Y(FE_PHN1684_key_mem_288_), 
	.A(key_mem[288]));
   DLY4X1 FE_PHC1683_key_mem_323_ (.Y(FE_PHN1683_key_mem_323_), 
	.A(key_mem[323]));
   DLY4X1 FE_PHC1682_key_mem_263_ (.Y(FE_PHN1682_key_mem_263_), 
	.A(key_mem[263]));
   DLY4X1 FE_PHC1681_n1552 (.Y(FE_PHN1681_n1552), 
	.A(FE_PHN4532_n1552));
   DLY4X1 FE_PHC1680_key_mem_734_ (.Y(FE_PHN1680_key_mem_734_), 
	.A(key_mem[734]));
   DLY4X1 FE_PHC1679_key_mem_757_ (.Y(FE_PHN1679_key_mem_757_), 
	.A(key_mem[757]));
   DLY4X1 FE_PHC1678_key_mem_715_ (.Y(FE_PHN1678_key_mem_715_), 
	.A(key_mem[715]));
   DLY4X1 FE_PHC1677_key_mem_363_ (.Y(FE_PHN1677_key_mem_363_), 
	.A(key_mem[363]));
   DLY4X1 FE_PHC1676_n1581 (.Y(FE_PHN1676_n1581), 
	.A(n1581));
   DLY4X1 FE_PHC1675_n1655 (.Y(FE_PHN1675_n1655), 
	.A(FE_PHN3871_n1655));
   DLY4X1 FE_PHC1674_n2172 (.Y(FE_PHN1674_n2172), 
	.A(FE_PHN4298_n2172));
   DLY4X1 FE_PHC1673_n1807 (.Y(FE_PHN1673_n1807), 
	.A(FE_PHN3890_n1807));
   DLY4X1 FE_PHC1672_key_mem_272_ (.Y(FE_PHN1672_key_mem_272_), 
	.A(key_mem[272]));
   DLY4X1 FE_PHC1671_key_mem_731_ (.Y(FE_PHN1671_key_mem_731_), 
	.A(key_mem[731]));
   DLY4X1 FE_PHC1670_key_mem_380_ (.Y(FE_PHN1670_key_mem_380_), 
	.A(key_mem[380]));
   DLY4X1 FE_PHC1669_n2077 (.Y(FE_PHN1669_n2077), 
	.A(FE_PHN3889_n2077));
   DLY4X1 FE_PHC1668_key_mem_742_ (.Y(FE_PHN1668_key_mem_742_), 
	.A(key_mem[742]));
   DLY4X1 FE_PHC1667_key_mem_322_ (.Y(FE_PHN1667_key_mem_322_), 
	.A(key_mem[322]));
   DLY4X1 FE_PHC1666_key_mem_730_ (.Y(FE_PHN1666_key_mem_730_), 
	.A(key_mem[730]));
   DLY4X1 FE_PHC1665_n2205 (.Y(FE_PHN1665_n2205), 
	.A(FE_PHN3876_n2205));
   DLY4X1 FE_PHC1664_n1461 (.Y(FE_PHN1664_n1461), 
	.A(FE_PHN4334_n1461));
   DLY4X1 FE_PHC1663_key_mem_687_ (.Y(FE_PHN1663_key_mem_687_), 
	.A(key_mem[687]));
   DLY4X1 FE_PHC1662_n1539 (.Y(FE_PHN1662_n1539), 
	.A(n1539));
   DLY4X1 FE_PHC1661_key_mem_677_ (.Y(FE_PHN1661_key_mem_677_), 
	.A(key_mem[677]));
   DLY4X1 FE_PHC1660_key_mem_663_ (.Y(FE_PHN1660_key_mem_663_), 
	.A(key_mem[663]));
   DLY4X1 FE_PHC1659_key_mem_354_ (.Y(FE_PHN1659_key_mem_354_), 
	.A(key_mem[354]));
   DLY4X1 FE_PHC1658_key_mem_317_ (.Y(FE_PHN1658_key_mem_317_), 
	.A(key_mem[317]));
   DLY4X1 FE_PHC1657_key_mem_656_ (.Y(FE_PHN1657_key_mem_656_), 
	.A(key_mem[656]));
   DLY4X1 FE_PHC1656_key_mem_701_ (.Y(FE_PHN1656_key_mem_701_), 
	.A(key_mem[701]));
   DLY4X1 FE_PHC1655_key_mem_358_ (.Y(FE_PHN1655_key_mem_358_), 
	.A(key_mem[358]));
   DLY4X1 FE_PHC1654_n1531 (.Y(FE_PHN1654_n1531), 
	.A(n1531));
   DLY4X1 FE_PHC1653_key_mem_342_ (.Y(FE_PHN1653_key_mem_342_), 
	.A(key_mem[342]));
   DLY4X1 FE_PHC1652_key_mem_261_ (.Y(FE_PHN1652_key_mem_261_), 
	.A(key_mem[261]));
   DLY4X1 FE_PHC1651_n2169 (.Y(FE_PHN1651_n2169), 
	.A(FE_PHN3848_n2169));
   DLY4X1 FE_PHC1650_key_mem_301_ (.Y(FE_PHN1650_key_mem_301_), 
	.A(key_mem[301]));
   DLY4X1 FE_PHC1649_n1671 (.Y(FE_PHN1649_n1671), 
	.A(FE_PHN3760_n1671));
   DLY4X1 FE_PHC1648_n2280 (.Y(FE_PHN1648_n2280), 
	.A(FE_PHN4242_n2280));
   DLY4X1 FE_PHC1647_n1520 (.Y(FE_PHN1647_n1520), 
	.A(FE_PHN4194_n1520));
   DLY4X1 FE_PHC1646_key_mem_726_ (.Y(FE_PHN1646_key_mem_726_), 
	.A(key_mem[726]));
   DLY4X1 FE_PHC1645_key_mem_697_ (.Y(FE_PHN1645_key_mem_697_), 
	.A(key_mem[697]));
   DLY4X1 FE_PHC1644_key_mem_370_ (.Y(FE_PHN1644_key_mem_370_), 
	.A(key_mem[370]));
   DLY4X1 FE_PHC1643_n1675 (.Y(FE_PHN1643_n1675), 
	.A(FE_PHN4355_n1675));
   DLY4X1 FE_PHC1642_key_mem_728_ (.Y(FE_PHN1642_key_mem_728_), 
	.A(key_mem[728]));
   DLY4X1 FE_PHC1641_key_mem_674_ (.Y(FE_PHN1641_key_mem_674_), 
	.A(key_mem[674]));
   DLY4X1 FE_PHC1640_n1745 (.Y(FE_PHN1640_n1745), 
	.A(FE_PHN3817_n1745));
   DLY4X1 FE_PHC1639_key_mem_274_ (.Y(FE_PHN1639_key_mem_274_), 
	.A(key_mem[274]));
   DLY4X1 FE_PHC1638_key_mem_692_ (.Y(FE_PHN1638_key_mem_692_), 
	.A(key_mem[692]));
   DLY4X1 FE_PHC1637_key_mem_338_ (.Y(FE_PHN1637_key_mem_338_), 
	.A(key_mem[338]));
   DLY4X1 FE_PHC1636_key_mem_750_ (.Y(FE_PHN1636_key_mem_750_), 
	.A(key_mem[750]));
   DLY4X1 FE_PHC1635_key_mem_315_ (.Y(FE_PHN1635_key_mem_315_), 
	.A(key_mem[315]));
   DLY4X1 FE_PHC1634_key_mem_280_ (.Y(FE_PHN1634_key_mem_280_), 
	.A(key_mem[280]));
   DLY4X1 FE_PHC1633_key_mem_307_ (.Y(FE_PHN1633_key_mem_307_), 
	.A(key_mem[307]));
   DLY4X1 FE_PHC1632_key_mem_264_ (.Y(FE_PHN1632_key_mem_264_), 
	.A(key_mem[264]));
   DLY4X1 FE_PHC1631_key_mem_756_ (.Y(FE_PHN1631_key_mem_756_), 
	.A(key_mem[756]));
   DLY4X1 FE_PHC1630_key_mem_685_ (.Y(FE_PHN1630_key_mem_685_), 
	.A(key_mem[685]));
   DLY4X1 FE_PHC1629_n2151 (.Y(FE_PHN1629_n2151), 
	.A(FE_PHN4203_n2151));
   DLY4X1 FE_PHC1628_n2125 (.Y(FE_PHN1628_n2125), 
	.A(n2125));
   DLY4X1 FE_PHC1627_key_mem_329_ (.Y(FE_PHN1627_key_mem_329_), 
	.A(key_mem[329]));
   DLY4X1 FE_PHC1626_key_mem_270_ (.Y(FE_PHN1626_key_mem_270_), 
	.A(key_mem[270]));
   DLY4X1 FE_PHC1625_n1618 (.Y(FE_PHN1625_n1618), 
	.A(FE_PHN3825_n1618));
   DLY4X1 FE_PHC1624_key_mem_645_ (.Y(FE_PHN1624_key_mem_645_), 
	.A(key_mem[645]));
   DLY4X1 FE_PHC1623_key_mem_281_ (.Y(FE_PHN1623_key_mem_281_), 
	.A(key_mem[281]));
   DLY4X1 FE_PHC1622_key_mem_278_ (.Y(FE_PHN1622_key_mem_278_), 
	.A(key_mem[278]));
   DLY4X1 FE_PHC1621_key_mem_321_ (.Y(FE_PHN1621_key_mem_321_), 
	.A(key_mem[321]));
   DLY4X1 FE_PHC1620_key_mem_340_ (.Y(FE_PHN1620_key_mem_340_), 
	.A(key_mem[340]));
   DLY4X1 FE_PHC1619_key_mem_355_ (.Y(FE_PHN1619_key_mem_355_), 
	.A(key_mem[355]));
   DLY4X1 FE_PHC1618_key_mem_365_ (.Y(FE_PHN1618_key_mem_365_), 
	.A(key_mem[365]));
   DLY4X1 FE_PHC1617_n2133 (.Y(FE_PHN1617_n2133), 
	.A(n2133));
   DLY4X1 FE_PHC1616_key_mem_293_ (.Y(FE_PHN1616_key_mem_293_), 
	.A(key_mem[293]));
   DLY4X1 FE_PHC1615_key_mem_643_ (.Y(FE_PHN1615_key_mem_643_), 
	.A(key_mem[643]));
   DLY4X1 FE_PHC1614_key_mem_350_ (.Y(FE_PHN1614_key_mem_350_), 
	.A(key_mem[350]));
   DLY4X1 FE_PHC1613_key_mem_751_ (.Y(FE_PHN1613_key_mem_751_), 
	.A(key_mem[751]));
   DLY4X1 FE_PHC1612_n2058 (.Y(FE_PHN1612_n2058), 
	.A(n2058));
   DLY4X1 FE_PHC1611_n1580 (.Y(FE_PHN1611_n1580), 
	.A(FE_PHN3933_n1580));
   DLY4X1 FE_PHC1610_n1908 (.Y(FE_PHN1610_n1908), 
	.A(FE_PHN4354_n1908));
   DLY4X1 FE_PHC1609_key_mem_711_ (.Y(FE_PHN1609_key_mem_711_), 
	.A(key_mem[711]));
   DLY4X1 FE_PHC1608_n2170 (.Y(FE_PHN1608_n2170), 
	.A(FE_PHN3898_n2170));
   DLY4X1 FE_PHC1607_key_mem_364_ (.Y(FE_PHN1607_key_mem_364_), 
	.A(key_mem[364]));
   DLY4X1 FE_PHC1606_key_mem_741_ (.Y(FE_PHN1606_key_mem_741_), 
	.A(key_mem[741]));
   DLY4X1 FE_PHC1605_key_mem_369_ (.Y(FE_PHN1605_key_mem_369_), 
	.A(key_mem[369]));
   DLY4X1 FE_PHC1604_n1660 (.Y(FE_PHN1604_n1660), 
	.A(FE_PHN3776_n1660));
   DLY4X1 FE_PHC1603_key_mem_330_ (.Y(FE_PHN1603_key_mem_330_), 
	.A(key_mem[330]));
   DLY4X1 FE_PHC1602_key_mem_765_ (.Y(FE_PHN1602_key_mem_765_), 
	.A(key_mem[765]));
   DLY4X1 FE_PHC1601_key_mem_294_ (.Y(FE_PHN1601_key_mem_294_), 
	.A(key_mem[294]));
   DLY4X1 FE_PHC1600_key_mem_303_ (.Y(FE_PHN1600_key_mem_303_), 
	.A(key_mem[303]));
   DLY4X1 FE_PHC1599_n2171 (.Y(FE_PHN1599_n2171), 
	.A(FE_PHN3703_n2171));
   DLY4X1 FE_PHC1598_key_mem_375_ (.Y(FE_PHN1598_key_mem_375_), 
	.A(key_mem[375]));
   DLY4X1 FE_PHC1597_n1750 (.Y(FE_PHN1597_n1750), 
	.A(FE_PHN3789_n1750));
   DLY4X1 FE_PHC1596_key_mem_735_ (.Y(FE_PHN1596_key_mem_735_), 
	.A(key_mem[735]));
   DLY4X1 FE_PHC1595_key_mem_361_ (.Y(FE_PHN1595_key_mem_361_), 
	.A(key_mem[361]));
   DLY4X1 FE_PHC1594_key_mem_362_ (.Y(FE_PHN1594_key_mem_362_), 
	.A(key_mem[362]));
   DLY4X1 FE_PHC1593_key_mem_686_ (.Y(FE_PHN1593_key_mem_686_), 
	.A(key_mem[686]));
   DLY4X1 FE_PHC1592_n1657 (.Y(FE_PHN1592_n1657), 
	.A(FE_PHN3784_n1657));
   DLY4X1 FE_PHC1591_n2064 (.Y(FE_PHN1591_n2064), 
	.A(FE_PHN4155_n2064));
   DLY4X1 FE_PHC1590_key_mem_752_ (.Y(FE_PHN1590_key_mem_752_), 
	.A(key_mem[752]));
   DLY4X1 FE_PHC1589_key_mem_378_ (.Y(FE_PHN1589_key_mem_378_), 
	.A(key_mem[378]));
   DLY4X1 FE_PHC1588_key_mem_655_ (.Y(FE_PHN1588_key_mem_655_), 
	.A(key_mem[655]));
   DLY4X1 FE_PHC1587_key_mem_733_ (.Y(FE_PHN1587_key_mem_733_), 
	.A(key_mem[733]));
   DLY4X1 FE_PHC1586_key_mem_298_ (.Y(FE_PHN1586_key_mem_298_), 
	.A(key_mem[298]));
   DLY4X1 FE_PHC1585_n1593 (.Y(FE_PHN1585_n1593), 
	.A(FE_PHN3830_n1593));
   DLY4X1 FE_PHC1584_key_mem_313_ (.Y(FE_PHN1584_key_mem_313_), 
	.A(key_mem[313]));
   DLY4X1 FE_PHC1583_key_mem_357_ (.Y(FE_PHN1583_key_mem_357_), 
	.A(key_mem[357]));
   DLY4X1 FE_PHC1582_n1545 (.Y(FE_PHN1582_n1545), 
	.A(FE_PHN4152_n1545));
   DLY4X1 FE_PHC1581_key_mem_672_ (.Y(FE_PHN1581_key_mem_672_), 
	.A(key_mem[672]));
   DLY4X1 FE_PHC1580_key_mem_372_ (.Y(FE_PHN1580_key_mem_372_), 
	.A(key_mem[372]));
   DLY4X1 FE_PHC1579_key_mem_678_ (.Y(FE_PHN1579_key_mem_678_), 
	.A(key_mem[678]));
   DLY4X1 FE_PHC1578_n1418 (.Y(FE_PHN1578_n1418), 
	.A(FE_PHN4186_n1418));
   DLY4X1 FE_PHC1577_key_mem_654_ (.Y(FE_PHN1577_key_mem_654_), 
	.A(key_mem[654]));
   DLY4X1 FE_PHC1576_n1546 (.Y(FE_PHN1576_n1546), 
	.A(n1546));
   DLY4X1 FE_PHC1575_key_mem_683_ (.Y(FE_PHN1575_key_mem_683_), 
	.A(key_mem[683]));
   DLY4X1 FE_PHC1574_key_mem_705_ (.Y(FE_PHN1574_key_mem_705_), 
	.A(key_mem[705]));
   DLY4X1 FE_PHC1573_key_mem_290_ (.Y(FE_PHN1573_key_mem_290_), 
	.A(key_mem[290]));
   DLY4X1 FE_PHC1572_key_mem_347_ (.Y(FE_PHN1572_key_mem_347_), 
	.A(key_mem[347]));
   DLY4X1 FE_PHC1571_key_mem_268_ (.Y(FE_PHN1571_key_mem_268_), 
	.A(key_mem[268]));
   DLY4X1 FE_PHC1570_n1577 (.Y(FE_PHN1570_n1577), 
	.A(FE_PHN3829_n1577));
   DLY4X1 FE_PHC1569_key_mem_670_ (.Y(FE_PHN1569_key_mem_670_), 
	.A(key_mem[670]));
   DLY4X1 FE_PHC1568_key_mem_720_ (.Y(FE_PHN1568_key_mem_720_), 
	.A(key_mem[720]));
   DLY4X1 FE_PHC1567_n2057 (.Y(FE_PHN1567_n2057), 
	.A(FE_PHN3678_n2057));
   DLY4X1 FE_PHC1566_n2264 (.Y(FE_PHN1566_n2264), 
	.A(FE_PHN3736_n2264));
   DLY4X1 FE_PHC1565_key_mem_679_ (.Y(FE_PHN1565_key_mem_679_), 
	.A(key_mem[679]));
   DLY4X1 FE_PHC1564_key_mem_681_ (.Y(FE_PHN1564_key_mem_681_), 
	.A(key_mem[681]));
   DLY4X1 FE_PHC1563_key_mem_368_ (.Y(FE_PHN1563_key_mem_368_), 
	.A(key_mem[368]));
   DLY4X1 FE_PHC1562_key_mem_296_ (.Y(FE_PHN1562_key_mem_296_), 
	.A(key_mem[296]));
   DLY4X1 FE_PHC1561_key_mem_706_ (.Y(FE_PHN1561_key_mem_706_), 
	.A(key_mem[706]));
   DLY4X1 FE_PHC1560_key_mem_811_ (.Y(FE_PHN1560_key_mem_811_), 
	.A(key_mem[811]));
   DLY4X1 FE_PHC1559_key_mem_306_ (.Y(FE_PHN1559_key_mem_306_), 
	.A(key_mem[306]));
   DLY4X1 FE_PHC1558_n2265 (.Y(FE_PHN1558_n2265), 
	.A(FE_PHN3811_n2265));
   DLY4X1 FE_PHC1557_key_mem_305_ (.Y(FE_PHN1557_key_mem_305_), 
	.A(key_mem[305]));
   DLY4X1 FE_PHC1556_key_mem_725_ (.Y(FE_PHN1556_key_mem_725_), 
	.A(key_mem[725]));
   DLY4X1 FE_PHC1555_key_mem_320_ (.Y(FE_PHN1555_key_mem_320_), 
	.A(key_mem[320]));
   DLY4X1 FE_PHC1554_key_mem_282_ (.Y(FE_PHN1554_key_mem_282_), 
	.A(key_mem[282]));
   DLY4X1 FE_PHC1553_key_mem_257_ (.Y(FE_PHN1553_key_mem_257_), 
	.A(key_mem[257]));
   DLY4X1 FE_PHC1552_key_mem_763_ (.Y(FE_PHN1552_key_mem_763_), 
	.A(key_mem[763]));
   DLY4X1 FE_PHC1551_n1739 (.Y(FE_PHN1551_n1739), 
	.A(FE_PHN3934_n1739));
   DLY4X1 FE_PHC1550_key_mem_744_ (.Y(FE_PHN1550_key_mem_744_), 
	.A(key_mem[744]));
   DLY4X1 FE_PHC1549_key_mem_356_ (.Y(FE_PHN1549_key_mem_356_), 
	.A(key_mem[356]));
   DLY4X1 FE_PHC1548_n2187 (.Y(FE_PHN1548_n2187), 
	.A(FE_PHN3730_n2187));
   DLY4X1 FE_PHC1547_key_mem_310_ (.Y(FE_PHN1547_key_mem_310_), 
	.A(key_mem[310]));
   DLY4X1 FE_PHC1546_key_mem_259_ (.Y(FE_PHN1546_key_mem_259_), 
	.A(key_mem[259]));
   DLY4X1 FE_PHC1545_key_mem_299_ (.Y(FE_PHN1545_key_mem_299_), 
	.A(key_mem[299]));
   DLY4X1 FE_PHC1544_key_mem_300_ (.Y(FE_PHN1544_key_mem_300_), 
	.A(key_mem[300]));
   DLY4X1 FE_PHC1543_key_mem_327_ (.Y(FE_PHN1543_key_mem_327_), 
	.A(key_mem[327]));
   DLY4X1 FE_PHC1542_key_mem_273_ (.Y(FE_PHN1542_key_mem_273_), 
	.A(key_mem[273]));
   DLY4X1 FE_PHC1541_n1447 (.Y(FE_PHN1541_n1447), 
	.A(n1447));
   DLY4X1 FE_PHC1540_n1419 (.Y(FE_PHN1540_n1419), 
	.A(FE_PHN4669_n1419));
   DLY4X1 FE_PHC1539_n1800 (.Y(FE_PHN1539_n1800), 
	.A(n1800));
   DLY4X1 FE_PHC1538_key_mem_366_ (.Y(FE_PHN1538_key_mem_366_), 
	.A(key_mem[366]));
   DLY4X1 FE_PHC1537_key_mem_312_ (.Y(FE_PHN1537_key_mem_312_), 
	.A(key_mem[312]));
   DLY4X1 FE_PHC1536_key_mem_754_ (.Y(FE_PHN1536_key_mem_754_), 
	.A(key_mem[754]));
   DLY4X1 FE_PHC1535_key_mem_699_ (.Y(FE_PHN1535_key_mem_699_), 
	.A(key_mem[699]));
   DLY4X1 FE_PHC1534_n1659 (.Y(FE_PHN1534_n1659), 
	.A(FE_PHN4084_n1659));
   DLY4X1 FE_PHC1533_key_mem_337_ (.Y(FE_PHN1533_key_mem_337_), 
	.A(key_mem[337]));
   DLY4X1 FE_PHC1532_key_mem_806_ (.Y(FE_PHN1532_key_mem_806_), 
	.A(key_mem[806]));
   DLY4X1 FE_PHC1531_key_mem_762_ (.Y(FE_PHN1531_key_mem_762_), 
	.A(key_mem[762]));
   DLY4X1 FE_PHC1530_key_mem_719_ (.Y(FE_PHN1530_key_mem_719_), 
	.A(key_mem[719]));
   DLY4X1 FE_PHC1529_key_mem_314_ (.Y(FE_PHN1529_key_mem_314_), 
	.A(key_mem[314]));
   DLY4X1 FE_PHC1528_key_mem_729_ (.Y(FE_PHN1528_key_mem_729_), 
	.A(key_mem[729]));
   DLY4X1 FE_PHC1527_n2183 (.Y(FE_PHN1527_n2183), 
	.A(FE_PHN3954_n2183));
   DLY4X1 FE_PHC1526_n2281 (.Y(FE_PHN1526_n2281), 
	.A(FE_PHN4022_n2281));
   DLY4X1 FE_PHC1525_key_mem_292_ (.Y(FE_PHN1525_key_mem_292_), 
	.A(key_mem[292]));
   DLY4X1 FE_PHC1524_key_mem_712_ (.Y(FE_PHN1524_key_mem_712_), 
	.A(key_mem[712]));
   DLY4X1 FE_PHC1523_key_mem_717_ (.Y(FE_PHN1523_key_mem_717_), 
	.A(key_mem[717]));
   DLY4X1 FE_PHC1522_key_mem_276_ (.Y(FE_PHN1522_key_mem_276_), 
	.A(key_mem[276]));
   DLY4X1 FE_PHC1521_key_mem_718_ (.Y(FE_PHN1521_key_mem_718_), 
	.A(key_mem[718]));
   DLY4X1 FE_PHC1520_key_mem_736_ (.Y(FE_PHN1520_key_mem_736_), 
	.A(key_mem[736]));
   DLY4X1 FE_PHC1519_key_mem_722_ (.Y(FE_PHN1519_key_mem_722_), 
	.A(key_mem[722]));
   DLY4X1 FE_PHC1518_key_mem_283_ (.Y(FE_PHN1518_key_mem_283_), 
	.A(key_mem[283]));
   DLY4X1 FE_PHC1517_key_mem_383_ (.Y(FE_PHN1517_key_mem_383_), 
	.A(key_mem[383]));
   DLY4X1 FE_PHC1516_key_mem_702_ (.Y(FE_PHN1516_key_mem_702_), 
	.A(key_mem[702]));
   DLY4X1 FE_PHC1515_key_mem_377_ (.Y(FE_PHN1515_key_mem_377_), 
	.A(key_mem[377]));
   DLY4X1 FE_PHC1514_key_mem_332_ (.Y(FE_PHN1514_key_mem_332_), 
	.A(key_mem[332]));
   DLY4X1 FE_PHC1513_n2048 (.Y(FE_PHN1513_n2048), 
	.A(FE_PHN4004_n2048));
   DLY4X1 FE_PHC1512_key_mem_664_ (.Y(FE_PHN1512_key_mem_664_), 
	.A(key_mem[664]));
   DLY4X1 FE_PHC1511_key_mem_295_ (.Y(FE_PHN1511_key_mem_295_), 
	.A(key_mem[295]));
   DLY4X1 FE_PHC1510_n1738 (.Y(FE_PHN1510_n1738), 
	.A(FE_PHN3864_n1738));
   DLY4X1 FE_PHC1509_n2147 (.Y(FE_PHN1509_n2147), 
	.A(FE_PHN4140_n2147));
   DLY4X1 FE_PHC1508_n1413 (.Y(FE_PHN1508_n1413), 
	.A(n1413));
   DLY4X1 FE_PHC1507_key_mem_304_ (.Y(FE_PHN1507_key_mem_304_), 
	.A(key_mem[304]));
   DLY4X1 FE_PHC1506_key_mem_690_ (.Y(FE_PHN1506_key_mem_690_), 
	.A(key_mem[690]));
   DLY4X1 FE_PHC1505_key_mem_658_ (.Y(FE_PHN1505_key_mem_658_), 
	.A(key_mem[658]));
   DLY4X1 FE_PHC1504_key_mem_271_ (.Y(FE_PHN1504_key_mem_271_), 
	.A(key_mem[271]));
   DLY4X1 FE_PHC1503_key_mem_382_ (.Y(FE_PHN1503_key_mem_382_), 
	.A(key_mem[382]));
   DLY4X1 FE_PHC1502_key_mem_642_ (.Y(FE_PHN1502_key_mem_642_), 
	.A(key_mem[642]));
   DLY4X1 FE_PHC1501_key_mem_381_ (.Y(FE_PHN1501_key_mem_381_), 
	.A(key_mem[381]));
   DLY4X1 FE_PHC1500_key_mem_749_ (.Y(FE_PHN1500_key_mem_749_), 
	.A(key_mem[749]));
   DLY4X1 FE_PHC1499_n2107 (.Y(FE_PHN1499_n2107), 
	.A(FE_PHN3700_n2107));
   DLY4X1 FE_PHC1498_key_mem_373_ (.Y(FE_PHN1498_key_mem_373_), 
	.A(key_mem[373]));
   DLY4X1 FE_PHC1497_n2042 (.Y(FE_PHN1497_n2042), 
	.A(FE_PHN3653_n2042));
   DLY4X1 FE_PHC1496_key_mem_319_ (.Y(FE_PHN1496_key_mem_319_), 
	.A(key_mem[319]));
   DLY4X1 FE_PHC1495_key_mem_714_ (.Y(FE_PHN1495_key_mem_714_), 
	.A(key_mem[714]));
   DLY4X1 FE_PHC1494_key_mem_335_ (.Y(FE_PHN1494_key_mem_335_), 
	.A(key_mem[335]));
   DLY4X1 FE_PHC1493_key_mem_336_ (.Y(FE_PHN1493_key_mem_336_), 
	.A(key_mem[336]));
   DLY4X1 FE_PHC1492_key_mem_289_ (.Y(FE_PHN1492_key_mem_289_), 
	.A(key_mem[289]));
   DLY4X1 FE_PHC1491_key_mem_840_ (.Y(FE_PHN1491_key_mem_840_), 
	.A(key_mem[840]));
   DLY4X1 FE_PHC1490_n2076 (.Y(FE_PHN1490_n2076), 
	.A(FE_PHN3657_n2076));
   DLY4X1 FE_PHC1489_n2263 (.Y(FE_PHN1489_n2263), 
	.A(FE_PHN3693_n2263));
   DLY4X1 FE_PHC1488_n2144 (.Y(FE_PHN1488_n2144), 
	.A(FE_PHN4196_n2144));
   DLY4X1 FE_PHC1487_n1667 (.Y(FE_PHN1487_n1667), 
	.A(FE_PHN3692_n1667));
   DLY4X1 FE_PHC1486_n1752 (.Y(FE_PHN1486_n1752), 
	.A(FE_PHN3720_n1752));
   DLY4X1 FE_PHC1485_n2063 (.Y(FE_PHN1485_n2063), 
	.A(FE_PHN4049_n2063));
   DLY4X1 FE_PHC1484_key_mem_277_ (.Y(FE_PHN1484_key_mem_277_), 
	.A(key_mem[277]));
   DLY4X1 FE_PHC1483_key_mem_700_ (.Y(FE_PHN1483_key_mem_700_), 
	.A(key_mem[700]));
   DLY4X1 FE_PHC1482_key_mem_284_ (.Y(FE_PHN1482_key_mem_284_), 
	.A(key_mem[284]));
   DLY4X1 FE_PHC1481_key_mem_649_ (.Y(FE_PHN1481_key_mem_649_), 
	.A(key_mem[649]));
   DLY4X1 FE_PHC1480_n1902 (.Y(FE_PHN1480_n1902), 
	.A(n1902));
   DLY4X1 FE_PHC1479_key_mem_326_ (.Y(FE_PHN1479_key_mem_326_), 
	.A(key_mem[326]));
   DLY4X1 FE_PHC1478_n2106 (.Y(FE_PHN1478_n2106), 
	.A(FE_PHN3702_n2106));
   DLY4X1 FE_PHC1477_key_mem_286_ (.Y(FE_PHN1477_key_mem_286_), 
	.A(key_mem[286]));
   DLY4X1 FE_PHC1476_key_mem_691_ (.Y(FE_PHN1476_key_mem_691_), 
	.A(key_mem[691]));
   DLY4X1 FE_PHC1475_key_mem_331_ (.Y(FE_PHN1475_key_mem_331_), 
	.A(key_mem[331]));
   DLY4X1 FE_PHC1474_n1737 (.Y(FE_PHN1474_n1737), 
	.A(FE_PHN3699_n1737));
   DLY4X1 FE_PHC1473_key_mem_748_ (.Y(FE_PHN1473_key_mem_748_), 
	.A(key_mem[748]));
   DLY4X1 FE_PHC1472_key_mem_333_ (.Y(FE_PHN1472_key_mem_333_), 
	.A(key_mem[333]));
   DLY4X1 FE_PHC1471_n2056 (.Y(FE_PHN1471_n2056), 
	.A(FE_PHN3658_n2056));
   DLY4X1 FE_PHC1470_n2050 (.Y(FE_PHN1470_n2050), 
	.A(FE_PHN3670_n2050));
   DLY4X1 FE_PHC1469_key_mem_835_ (.Y(FE_PHN1469_key_mem_835_), 
	.A(key_mem[835]));
   DLY4X1 FE_PHC1468_n2266 (.Y(FE_PHN1468_n2266), 
	.A(FE_PHN3624_n2266));
   DLY4X1 FE_PHC1467_n1658 (.Y(FE_PHN1467_n1658), 
	.A(FE_PHN3620_n1658));
   DLY4X1 FE_PHC1466_n2124 (.Y(FE_PHN1466_n2124), 
	.A(FE_PHN3639_n2124));
   DLY4X1 FE_PHC1464_key_mem_339_ (.Y(FE_PHN1464_key_mem_339_), 
	.A(key_mem[339]));
   DLY4X1 FE_PHC1463_n2399 (.Y(FE_PHN1463_n2399), 
	.A(FE_PHN5057_n2399));
   DLY4X1 FE_PHC1446_prev_key1_reg_68_ (.Y(FE_PHN1446_prev_key1_reg_68_), 
	.A(prev_key1_reg[68]));
   DLY4X1 FE_PHC1445_prev_key1_reg_69_ (.Y(FE_PHN1445_prev_key1_reg_69_), 
	.A(prev_key1_reg[69]));
   DLY4X1 FE_PHC1444_prev_key1_reg_67_ (.Y(FE_PHN1444_prev_key1_reg_67_), 
	.A(prev_key1_reg[67]));
   DLY4X1 FE_PHC1442_prev_key1_reg_66_ (.Y(FE_PHN1442_prev_key1_reg_66_), 
	.A(prev_key1_reg[66]));
   DLY4X1 FE_PHC1441_prev_key1_reg_64_ (.Y(FE_PHN1441_prev_key1_reg_64_), 
	.A(prev_key1_reg[64]));
   DLY4X1 FE_PHC1434_prev_key1_reg_127_ (.Y(FE_PHN1434_prev_key1_reg_127_), 
	.A(prev_key1_reg[127]));
   DLY4X1 FE_PHC1429_prev_key1_reg_76_ (.Y(FE_PHN1429_prev_key1_reg_76_), 
	.A(prev_key1_reg[76]));
   DLY4X1 FE_PHC1425_prev_key1_reg_81_ (.Y(FE_PHN1425_prev_key1_reg_81_), 
	.A(prev_key1_reg[81]));
   DLY4X1 FE_PHC1421_prev_key1_reg_124_ (.Y(FE_PHN1421_prev_key1_reg_124_), 
	.A(prev_key1_reg[124]));
   DLY4X1 FE_PHC1416_prev_key1_reg_120_ (.Y(FE_PHN1416_prev_key1_reg_120_), 
	.A(prev_key1_reg[120]));
   DLY4X1 FE_PHC1415_prev_key1_reg_75_ (.Y(FE_PHN1415_prev_key1_reg_75_), 
	.A(prev_key1_reg[75]));
   DLY4X1 FE_PHC1414_prev_key1_reg_80_ (.Y(FE_PHN1414_prev_key1_reg_80_), 
	.A(prev_key1_reg[80]));
   DLY4X1 FE_PHC1413_prev_key1_reg_123_ (.Y(FE_PHN1413_prev_key1_reg_123_), 
	.A(prev_key1_reg[123]));
   DLY4X1 FE_PHC1412_prev_key1_reg_85_ (.Y(FE_PHN1412_prev_key1_reg_85_), 
	.A(prev_key1_reg[85]));
   DLY4X1 FE_PHC1408_prev_key1_reg_74_ (.Y(FE_PHN1408_prev_key1_reg_74_), 
	.A(prev_key1_reg[74]));
   DLY4X1 FE_PHC1406_prev_key1_reg_71_ (.Y(FE_PHN1406_prev_key1_reg_71_), 
	.A(prev_key1_reg[71]));
   DLY4X1 FE_PHC1405_prev_key1_reg_82_ (.Y(FE_PHN1405_prev_key1_reg_82_), 
	.A(prev_key1_reg[82]));
   DLY4X1 FE_PHC1404_prev_key1_reg_72_ (.Y(FE_PHN1404_prev_key1_reg_72_), 
	.A(prev_key1_reg[72]));
   DLY4X1 FE_PHC1402_prev_key1_reg_78_ (.Y(FE_PHN1402_prev_key1_reg_78_), 
	.A(prev_key1_reg[78]));
   DLY4X1 FE_PHC1401_prev_key1_reg_73_ (.Y(FE_PHN1401_prev_key1_reg_73_), 
	.A(prev_key1_reg[73]));
   DLY4X1 FE_PHC1397_prev_key1_reg_77_ (.Y(FE_PHN1397_prev_key1_reg_77_), 
	.A(prev_key1_reg[77]));
   DLY4X1 FE_PHC1395_prev_key1_reg_121_ (.Y(FE_PHN1395_prev_key1_reg_121_), 
	.A(prev_key1_reg[121]));
   DLY4X1 FE_PHC1394_prev_key1_reg_65_ (.Y(FE_PHN1394_prev_key1_reg_65_), 
	.A(prev_key1_reg[65]));
   DLY4X1 FE_PHC1393_prev_key1_reg_79_ (.Y(FE_PHN1393_prev_key1_reg_79_), 
	.A(prev_key1_reg[79]));
   DLY4X1 FE_PHC1392_prev_key1_reg_122_ (.Y(FE_PHN1392_prev_key1_reg_122_), 
	.A(prev_key1_reg[122]));
   DLY4X1 FE_PHC1391_prev_key1_reg_125_ (.Y(FE_PHN1391_prev_key1_reg_125_), 
	.A(prev_key1_reg[125]));
   DLY4X1 FE_PHC1388_prev_key1_reg_83_ (.Y(FE_PHN1388_prev_key1_reg_83_), 
	.A(prev_key1_reg[83]));
   DLY4X1 FE_PHC1375_prev_key1_reg_84_ (.Y(FE_PHN1375_prev_key1_reg_84_), 
	.A(prev_key1_reg[84]));
   DLY4X1 FE_PHC1333_n1283 (.Y(FE_PHN1333_n1283), 
	.A(FE_PHN4713_n1283));
   DLY4X1 FE_PHC1326_n1227 (.Y(FE_PHN1326_n1227), 
	.A(FE_PHN4362_n1227));
   DLY4X1 FE_PHC1324_n1029 (.Y(FE_PHN1324_n1029), 
	.A(n1029));
   DLY4X1 FE_PHC1323_n1163 (.Y(FE_PHN1323_n1163), 
	.A(FE_PHN4508_n1163));
   DLY4X1 FE_PHC1322_n1030 (.Y(FE_PHN1322_n1030), 
	.A(n1030));
   DLY4X1 FE_PHC1321_n971 (.Y(FE_PHN1321_n971), 
	.A(FE_PHN4139_n971));
   DLY4X1 FE_PHC1318_n972 (.Y(FE_PHN1318_n972), 
	.A(FE_PHN3978_n972));
   DLY4X1 FE_PHC1315_n2373 (.Y(FE_PHN1315_n2373), 
	.A(n2373));
   DLY4X1 FE_PHC1314_prev_key1_reg_119_ (.Y(FE_PHN1314_prev_key1_reg_119_), 
	.A(prev_key1_reg[119]));
   DLY4X1 FE_PHC1313_prev_key1_reg_118_ (.Y(FE_PHN1313_prev_key1_reg_118_), 
	.A(prev_key1_reg[118]));
   DLY4X1 FE_PHC1312_n2381 (.Y(FE_PHN1312_n2381), 
	.A(n2381));
   DLY4X1 FE_PHC1311_n1967 (.Y(FE_PHN1311_n1967), 
	.A(FE_PHN3774_n1967));
   DLY4X1 FE_PHC1263_rcon_reg_1_ (.Y(FE_PHN1263_rcon_reg_1_), 
	.A(rcon_reg[1]));
   DLY4X1 FE_PHC1257_rcon_reg_4_ (.Y(FE_PHN1257_rcon_reg_4_), 
	.A(rcon_reg[4]));
   DLY4X1 FE_PHC1256_prev_key1_reg_112_ (.Y(FE_PHN1256_prev_key1_reg_112_), 
	.A(prev_key1_reg[112]));
   DLY4X1 FE_PHC1252_prev_key1_reg_105_ (.Y(FE_PHN1252_prev_key1_reg_105_), 
	.A(prev_key1_reg[105]));
   DLY4X1 FE_PHC1251_prev_key1_reg_108_ (.Y(FE_PHN1251_prev_key1_reg_108_), 
	.A(prev_key1_reg[108]));
   DLY4X1 FE_PHC1249_prev_key1_reg_116_ (.Y(FE_PHN1249_prev_key1_reg_116_), 
	.A(prev_key1_reg[116]));
   DLY4X1 FE_PHC1246_n1736 (.Y(FE_PHN1246_n1736), 
	.A(FE_PHN4064_n1736));
   DLY4X1 FE_PHC1245_prev_key1_reg_99_ (.Y(FE_PHN1245_prev_key1_reg_99_), 
	.A(prev_key1_reg[99]));
   DLY4X1 FE_PHC1244_prev_key1_reg_115_ (.Y(FE_PHN1244_prev_key1_reg_115_), 
	.A(prev_key1_reg[115]));
   DLY4X1 FE_PHC1241_rcon_reg_5_ (.Y(FE_PHN1241_rcon_reg_5_), 
	.A(rcon_reg[5]));
   DLY4X1 FE_PHC1239_prev_key1_reg_97_ (.Y(FE_PHN1239_prev_key1_reg_97_), 
	.A(prev_key1_reg[97]));
   DLY4X1 FE_PHC1238_prev_key1_reg_98_ (.Y(FE_PHN1238_prev_key1_reg_98_), 
	.A(prev_key1_reg[98]));
   DLY4X1 FE_PHC1236_prev_key1_reg_113_ (.Y(FE_PHN1236_prev_key1_reg_113_), 
	.A(prev_key1_reg[113]));
   DLY4X1 FE_PHC1235_prev_key1_reg_117_ (.Y(FE_PHN1235_prev_key1_reg_117_), 
	.A(prev_key1_reg[117]));
   DLY4X1 FE_PHC1234_prev_key1_reg_109_ (.Y(FE_PHN1234_prev_key1_reg_109_), 
	.A(prev_key1_reg[109]));
   DLY4X1 FE_PHC1233_prev_key1_reg_106_ (.Y(FE_PHN1233_prev_key1_reg_106_), 
	.A(prev_key1_reg[106]));
   DLY4X1 FE_PHC1232_prev_key1_reg_107_ (.Y(FE_PHN1232_prev_key1_reg_107_), 
	.A(prev_key1_reg[107]));
   DLY4X1 FE_PHC1231_prev_key1_reg_96_ (.Y(FE_PHN1231_prev_key1_reg_96_), 
	.A(prev_key1_reg[96]));
   DLY4X1 FE_PHC1230_prev_key1_reg_53_ (.Y(FE_PHN1230_prev_key1_reg_53_), 
	.A(prev_key1_reg[53]));
   DLY4X1 FE_PHC1229_prev_key1_reg_101_ (.Y(FE_PHN1229_prev_key1_reg_101_), 
	.A(prev_key1_reg[101]));
   DLY4X1 FE_PHC1227_n2279 (.Y(FE_PHN1227_n2279), 
	.A(FE_PHN4054_n2279));
   DLY4X1 FE_PHC1226_prev_key1_reg_114_ (.Y(FE_PHN1226_prev_key1_reg_114_), 
	.A(prev_key1_reg[114]));
   DLY4X1 FE_PHC1225_prev_key1_reg_100_ (.Y(FE_PHN1225_prev_key1_reg_100_), 
	.A(prev_key1_reg[100]));
   DLY4X1 FE_PHC1224_prev_key1_reg_103_ (.Y(FE_PHN1224_prev_key1_reg_103_), 
	.A(prev_key1_reg[103]));
   DLY4X1 FE_PHC1223_prev_key1_reg_104_ (.Y(FE_PHN1223_prev_key1_reg_104_), 
	.A(prev_key1_reg[104]));
   DLY4X1 FE_PHC1221_prev_key1_reg_111_ (.Y(FE_PHN1221_prev_key1_reg_111_), 
	.A(prev_key1_reg[111]));
   DLY4X1 FE_PHC1220_prev_key1_reg_102_ (.Y(FE_PHN1220_prev_key1_reg_102_), 
	.A(prev_key1_reg[102]));
   DLY4X1 FE_PHC1219_prev_key1_reg_110_ (.Y(FE_PHN1219_prev_key1_reg_110_), 
	.A(prev_key1_reg[110]));
   DLY4X1 FE_PHC1211_n2294 (.Y(FE_PHN1211_n2294), 
	.A(FE_PHN4993_n2294));
   DLY4X1 FE_PHC1164_n1282 (.Y(FE_PHN1164_n1282), 
	.A(FE_PHN4838_n1282));
   DLY4X1 FE_PHC1100_n1288 (.Y(FE_PHN1100_n1288), 
	.A(FE_PHN4383_n1288));
   DLY4X1 FE_PHC1098_n1170 (.Y(FE_PHN1098_n1170), 
	.A(FE_PHN4512_n1170));
   DLY4X1 FE_PHC1096_n1022 (.Y(FE_PHN1096_n1022), 
	.A(n1022));
   DLY4X1 FE_PHC1093_n1153 (.Y(FE_PHN1093_n1153), 
	.A(FE_PHN4506_n1153));
   DLY4X1 FE_PHC1092_n1296 (.Y(FE_PHN1092_n1296), 
	.A(FE_PHN4352_n1296));
   DLY4X1 FE_PHC1088_n1295 (.Y(FE_PHN1088_n1295), 
	.A(FE_PHN4431_n1295));
   DLY4X1 FE_PHC1087_prev_key1_reg_44_ (.Y(FE_PHN1087_prev_key1_reg_44_), 
	.A(prev_key1_reg[44]));
   DLY4X1 FE_PHC1086_n1166 (.Y(FE_PHN1086_n1166), 
	.A(FE_PHN4424_n1166));
   DLY4X1 FE_PHC1085_n1041 (.Y(FE_PHN1085_n1041), 
	.A(FE_PHN3928_n1041));
   DLY4X1 FE_PHC1084_n1013 (.Y(FE_PHN1084_n1013), 
	.A(n1013));
   DLY4X1 FE_PHC1083_key_mem_1189_ (.Y(FE_PHN1083_key_mem_1189_), 
	.A(key_mem[1189]));
   DLY4X1 FE_PHC1081_n1299 (.Y(FE_PHN1081_n1299), 
	.A(FE_PHN4145_n1299));
   DLY4X1 FE_PHC1080_n1280 (.Y(FE_PHN1080_n1280), 
	.A(FE_PHN4286_n1280));
   DLY4X1 FE_PHC1079_prev_key1_reg_32_ (.Y(FE_PHN1079_prev_key1_reg_32_), 
	.A(prev_key1_reg[32]));
   DLY4X1 FE_PHC1077_n991 (.Y(FE_PHN1077_n991), 
	.A(FE_PHN4057_n991));
   DLY4X1 FE_PHC1076_n1023 (.Y(FE_PHN1076_n1023), 
	.A(FE_PHN4040_n1023));
   DLY4X1 FE_PHC1075_n1290 (.Y(FE_PHN1075_n1290), 
	.A(n1290));
   DLY4X1 FE_PHC1074_prev_key1_reg_50_ (.Y(FE_PHN1074_prev_key1_reg_50_), 
	.A(prev_key1_reg[50]));
   DLY4X1 FE_PHC1067_prev_key1_reg_49_ (.Y(FE_PHN1067_prev_key1_reg_49_), 
	.A(prev_key1_reg[49]));
   DLY4X1 FE_PHC1066_n908 (.Y(FE_PHN1066_n908), 
	.A(FE_PHN3866_n908));
   DLY4X1 FE_PHC1064_prev_key1_reg_45_ (.Y(FE_PHN1064_prev_key1_reg_45_), 
	.A(prev_key1_reg[45]));
   DLY4X1 FE_PHC1063_prev_key1_reg_35_ (.Y(FE_PHN1063_prev_key1_reg_35_), 
	.A(prev_key1_reg[35]));
   DLY4X1 FE_PHC1062_prev_key1_reg_47_ (.Y(FE_PHN1062_prev_key1_reg_47_), 
	.A(prev_key1_reg[47]));
   DLY4X1 FE_PHC1060_prev_key1_reg_33_ (.Y(FE_PHN1060_prev_key1_reg_33_), 
	.A(prev_key1_reg[33]));
   DLY4X1 FE_PHC1058_prev_key1_reg_41_ (.Y(FE_PHN1058_prev_key1_reg_41_), 
	.A(prev_key1_reg[41]));
   DLY4X1 FE_PHC1057_prev_key1_reg_55_ (.Y(FE_PHN1057_prev_key1_reg_55_), 
	.A(prev_key1_reg[55]));
   DLY4X1 FE_PHC1056_prev_key1_reg_37_ (.Y(FE_PHN1056_prev_key1_reg_37_), 
	.A(prev_key1_reg[37]));
   DLY4X1 FE_PHC1055_prev_key1_reg_38_ (.Y(FE_PHN1055_prev_key1_reg_38_), 
	.A(prev_key1_reg[38]));
   DLY4X1 FE_PHC1054_prev_key1_reg_42_ (.Y(FE_PHN1054_prev_key1_reg_42_), 
	.A(prev_key1_reg[42]));
   DLY4X1 FE_PHC1053_prev_key1_reg_36_ (.Y(FE_PHN1053_prev_key1_reg_36_), 
	.A(prev_key1_reg[36]));
   DLY4X1 FE_PHC1052_prev_key1_reg_51_ (.Y(FE_PHN1052_prev_key1_reg_51_), 
	.A(prev_key1_reg[51]));
   DLY4X1 FE_PHC1051_prev_key1_reg_40_ (.Y(FE_PHN1051_prev_key1_reg_40_), 
	.A(prev_key1_reg[40]));
   DLY4X1 FE_PHC1050_prev_key1_reg_54_ (.Y(FE_PHN1050_prev_key1_reg_54_), 
	.A(prev_key1_reg[54]));
   DLY4X1 FE_PHC1049_prev_key1_reg_39_ (.Y(FE_PHN1049_prev_key1_reg_39_), 
	.A(prev_key1_reg[39]));
   DLY4X1 FE_PHC1048_prev_key1_reg_43_ (.Y(FE_PHN1048_prev_key1_reg_43_), 
	.A(prev_key1_reg[43]));
   DLY4X1 FE_PHC1046_n2061 (.Y(FE_PHN1046_n2061), 
	.A(FE_PHN4220_n2061));
   DLY4X1 FE_PHC1045_n1782 (.Y(FE_PHN1045_n1782), 
	.A(FE_PHN4107_n1782));
   DLY4X1 FE_PHC1044_prev_key1_reg_34_ (.Y(FE_PHN1044_prev_key1_reg_34_), 
	.A(prev_key1_reg[34]));
   DLY4X1 FE_PHC1043_prev_key1_reg_52_ (.Y(FE_PHN1043_prev_key1_reg_52_), 
	.A(prev_key1_reg[52]));
   DLY4X1 FE_PHC1041_n1808 (.Y(FE_PHN1041_n1808), 
	.A(FE_PHN4167_n1808));
   DLY4X1 FE_PHC1040_n1766 (.Y(FE_PHN1040_n1766), 
	.A(FE_PHN4198_n1766));
   DLY4X1 FE_PHC1038_n2418 (.Y(FE_PHN1038_n2418), 
	.A(FE_PHN5030_n2418));
   DLY4X1 FE_PHC1037_n2432 (.Y(FE_PHN1037_n2432), 
	.A(n2432));
   DLY4X1 FE_PHC1036_rcon_reg_3_ (.Y(FE_PHN1036_rcon_reg_3_), 
	.A(rcon_reg[3]));
   DLY4X1 FE_PHC1035_n2350 (.Y(FE_PHN1035_n2350), 
	.A(FE_PHN4984_n2350));
   DLY4X1 FE_PHC1034_rcon_reg_0_ (.Y(FE_PHN1034_rcon_reg_0_), 
	.A(rcon_reg[0]));
   DLY4X1 FE_PHC1033_rcon_reg_2_ (.Y(FE_PHN1033_rcon_reg_2_), 
	.A(rcon_reg[2]));
   DLY4X1 FE_PHC1032_n2868 (.Y(FE_PHN1032_n2868), 
	.A(FE_PHN3373_n2868));
   DLY4X1 FE_PHC1029_key_mem_1193_ (.Y(FE_PHN1029_key_mem_1193_), 
	.A(key_mem[1193]));
   DLY4X1 FE_PHC1024_key_mem_1205_ (.Y(FE_PHN1024_key_mem_1205_), 
	.A(key_mem[1205]));
   DLY4X1 FE_PHC1023_key_mem_1155_ (.Y(FE_PHN1023_key_mem_1155_), 
	.A(key_mem[1155]));
   DLY4X1 FE_PHC1022_n1268 (.Y(FE_PHN1022_n1268), 
	.A(FE_PHN4944_n1268));
   DLY4X1 FE_PHC1021_key_mem_1206_ (.Y(FE_PHN1021_key_mem_1206_), 
	.A(key_mem[1206]));
   DLY4X1 FE_PHC1016_n1201 (.Y(FE_PHN1016_n1201), 
	.A(FE_PHN4509_n1201));
   DLY4X1 FE_PHC1015_key_mem_1186_ (.Y(FE_PHN1015_key_mem_1186_), 
	.A(key_mem[1186]));
   DLY4X1 FE_PHC1014_key_mem_1253_ (.Y(FE_PHN1014_key_mem_1253_), 
	.A(key_mem[1253]));
   DLY4X1 FE_PHC1011_n1076 (.Y(FE_PHN1011_n1076), 
	.A(FE_PHN4439_n1076));
   DLY4X1 FE_PHC1010_key_mem_1222_ (.Y(FE_PHN1010_key_mem_1222_), 
	.A(key_mem[1222]));
   DLY4X1 FE_PHC1009_key_mem_1259_ (.Y(FE_PHN1009_key_mem_1259_), 
	.A(key_mem[1259]));
   DLY4X1 FE_PHC1008_key_mem_1199_ (.Y(FE_PHN1008_key_mem_1199_), 
	.A(key_mem[1199]));
   DLY4X1 FE_PHC1006_key_mem_1219_ (.Y(FE_PHN1006_key_mem_1219_), 
	.A(key_mem[1219]));
   DLY4X1 FE_PHC1005_key_mem_1192_ (.Y(FE_PHN1005_key_mem_1192_), 
	.A(key_mem[1192]));
   DLY4X1 FE_PHC1000_key_mem_1174_ (.Y(FE_PHN1000_key_mem_1174_), 
	.A(key_mem[1174]));
   DLY4X1 FE_PHC999_n1182 (.Y(FE_PHN999_n1182), 
	.A(FE_PHN4600_n1182));
   DLY4X1 FE_PHC998_n1376 (.Y(FE_PHN998_n1376), 
	.A(FE_PHN4493_n1376));
   DLY4X1 FE_PHC997_n1386 (.Y(FE_PHN997_n1386), 
	.A(FE_PHN4521_n1386));
   DLY4X1 FE_PHC996_n1265 (.Y(FE_PHN996_n1265), 
	.A(FE_PHN4391_n1265));
   DLY4X1 FE_PHC995_n1320 (.Y(FE_PHN995_n1320), 
	.A(FE_PHN4137_n1320));
   DLY4X1 FE_PHC994_n888 (.Y(FE_PHN994_n888), 
	.A(FE_PHN4128_n888));
   DLY4X1 FE_PHC993_n1379 (.Y(FE_PHN993_n1379), 
	.A(FE_PHN4515_n1379));
   DLY4X1 FE_PHC992_key_mem_1202_ (.Y(FE_PHN992_key_mem_1202_), 
	.A(key_mem[1202]));
   DLY4X1 FE_PHC991_n1306 (.Y(FE_PHN991_n1306), 
	.A(FE_PHN4356_n1306));
   DLY4X1 FE_PHC990_key_mem_1270_ (.Y(FE_PHN990_key_mem_1270_), 
	.A(key_mem[1270]));
   DLY4X1 FE_PHC989_key_mem_1157_ (.Y(FE_PHN989_key_mem_1157_), 
	.A(key_mem[1157]));
   DLY4X1 FE_PHC988_n1391 (.Y(FE_PHN988_n1391), 
	.A(FE_PHN4364_n1391));
   DLY4X1 FE_PHC986_n1121 (.Y(FE_PHN986_n1121), 
	.A(n1121));
   DLY4X1 FE_PHC984_key_mem_1271_ (.Y(FE_PHN984_key_mem_1271_), 
	.A(key_mem[1271]));
   DLY4X1 FE_PHC983_n1331 (.Y(FE_PHN983_n1331), 
	.A(FE_PHN4568_n1331));
   DLY4X1 FE_PHC982_n1017 (.Y(FE_PHN982_n1017), 
	.A(FE_PHN4246_n1017));
   DLY4X1 FE_PHC981_key_mem_1261_ (.Y(FE_PHN981_key_mem_1261_), 
	.A(key_mem[1261]));
   DLY4X1 FE_PHC980_key_mem_1158_ (.Y(FE_PHN980_key_mem_1158_), 
	.A(key_mem[1158]));
   DLY4X1 FE_PHC979_prev_key1_reg_88_ (.Y(FE_PHN979_prev_key1_reg_88_), 
	.A(prev_key1_reg[88]));
   DLY4X1 FE_PHC977_key_mem_1220_ (.Y(FE_PHN977_key_mem_1220_), 
	.A(key_mem[1220]));
   DLY4X1 FE_PHC976_n892 (.Y(FE_PHN976_n892), 
	.A(n892));
   DLY4X1 FE_PHC975_key_mem_1227_ (.Y(FE_PHN975_key_mem_1227_), 
	.A(key_mem[1227]));
   DLY4X1 FE_PHC974_key_mem_1163_ (.Y(FE_PHN974_key_mem_1163_), 
	.A(key_mem[1163]));
   DLY4X1 FE_PHC973_n1196 (.Y(FE_PHN973_n1196), 
	.A(FE_PHN4072_n1196));
   DLY4X1 FE_PHC972_key_mem_1235_ (.Y(FE_PHN972_key_mem_1235_), 
	.A(key_mem[1235]));
   DLY4X1 FE_PHC971_n1012 (.Y(FE_PHN971_n1012), 
	.A(FE_PHN4032_n1012));
   DLY4X1 FE_PHC970_n1055 (.Y(FE_PHN970_n1055), 
	.A(FE_PHN4052_n1055));
   DLY4X1 FE_PHC969_key_mem_1344_ (.Y(FE_PHN969_key_mem_1344_), 
	.A(key_mem[1344]));
   DLY4X1 FE_PHC968_key_mem_1236_ (.Y(FE_PHN968_key_mem_1236_), 
	.A(key_mem[1236]));
   DLY4X1 FE_PHC966_n1385 (.Y(FE_PHN966_n1385), 
	.A(FE_PHN4208_n1385));
   DLY4X1 FE_PHC965_key_mem_1266_ (.Y(FE_PHN965_key_mem_1266_), 
	.A(key_mem[1266]));
   DLY4X1 FE_PHC964_n1688 (.Y(FE_PHN964_n1688), 
	.A(FE_PHN4478_n1688));
   DLY4X1 FE_PHC963_n1124 (.Y(FE_PHN963_n1124), 
	.A(FE_PHN4164_n1124));
   DLY4X1 FE_PHC962_n1184 (.Y(FE_PHN962_n1184), 
	.A(FE_PHN4381_n1184));
   DLY4X1 FE_PHC961_n1143 (.Y(FE_PHN961_n1143), 
	.A(FE_PHN4010_n1143));
   DLY4X1 FE_PHC960_key_mem_1228_ (.Y(FE_PHN960_key_mem_1228_), 
	.A(key_mem[1228]));
   DLY4X1 FE_PHC959_n1254 (.Y(FE_PHN959_n1254), 
	.A(FE_PHN4115_n1254));
   DLY4X1 FE_PHC958_key_mem_1201_ (.Y(FE_PHN958_key_mem_1201_), 
	.A(key_mem[1201]));
   DLY4X1 FE_PHC957_n1396 (.Y(FE_PHN957_n1396), 
	.A(FE_PHN4318_n1396));
   DLY4X1 FE_PHC956_n1128 (.Y(FE_PHN956_n1128), 
	.A(FE_PHN4025_n1128));
   DLY4X1 FE_PHC955_key_mem_1198_ (.Y(FE_PHN955_key_mem_1198_), 
	.A(key_mem[1198]));
   DLY4X1 FE_PHC954_key_mem_1063_ (.Y(FE_PHN954_key_mem_1063_), 
	.A(key_mem[1063]));
   DLY4X1 FE_PHC953_key_mem_1200_ (.Y(FE_PHN953_key_mem_1200_), 
	.A(key_mem[1200]));
   DLY4X1 FE_PHC950_n891 (.Y(FE_PHN950_n891), 
	.A(n891));
   DLY4X1 FE_PHC949_key_mem_1231_ (.Y(FE_PHN949_key_mem_1231_), 
	.A(key_mem[1231]));
   DLY4X1 FE_PHC948_n1395 (.Y(FE_PHN948_n1395), 
	.A(FE_PHN4058_n1395));
   DLY4X1 FE_PHC947_key_mem_1260_ (.Y(FE_PHN947_key_mem_1260_), 
	.A(key_mem[1260]));
   DLY4X1 FE_PHC945_n1185 (.Y(FE_PHN945_n1185), 
	.A(FE_PHN4047_n1185));
   DLY4X1 FE_PHC944_n1127 (.Y(FE_PHN944_n1127), 
	.A(FE_PHN4116_n1127));
   DLY4X1 FE_PHC943_key_mem_1195_ (.Y(FE_PHN943_key_mem_1195_), 
	.A(key_mem[1195]));
   DLY4X1 FE_PHC942_key_mem_1203_ (.Y(FE_PHN942_key_mem_1203_), 
	.A(key_mem[1203]));
   DLY4X1 FE_PHC940_prev_key1_reg_95_ (.Y(FE_PHN940_prev_key1_reg_95_), 
	.A(prev_key1_reg[95]));
   DLY4X1 FE_PHC939_key_mem_695_ (.Y(FE_PHN939_key_mem_695_), 
	.A(key_mem[695]));
   DLY4X1 FE_PHC938_n944 (.Y(FE_PHN938_n944), 
	.A(FE_PHN4018_n944));
   DLY4X1 FE_PHC937_n990 (.Y(FE_PHN937_n990), 
	.A(n990));
   DLY4X1 FE_PHC936_key_mem_1238_ (.Y(FE_PHN936_key_mem_1238_), 
	.A(key_mem[1238]));
   DLY4X1 FE_PHC935_key_mem_1268_ (.Y(FE_PHN935_key_mem_1268_), 
	.A(key_mem[1268]));
   DLY4X1 FE_PHC934_key_mem_1229_ (.Y(FE_PHN934_key_mem_1229_), 
	.A(key_mem[1229]));
   DLY4X1 FE_PHC933_prev_key1_reg_94_ (.Y(FE_PHN933_prev_key1_reg_94_), 
	.A(prev_key1_reg[94]));
   DLY4X1 FE_PHC932_key_mem_1379_ (.Y(FE_PHN932_key_mem_1379_), 
	.A(key_mem[1379]));
   DLY4X1 FE_PHC930_n946 (.Y(FE_PHN930_n946), 
	.A(FE_PHN3986_n946));
   DLY4X1 FE_PHC929_key_mem_1196_ (.Y(FE_PHN929_key_mem_1196_), 
	.A(key_mem[1196]));
   DLY4X1 FE_PHC928_n994 (.Y(FE_PHN928_n994), 
	.A(n994));
   DLY4X1 FE_PHC924_prev_key1_reg_90_ (.Y(FE_PHN924_prev_key1_reg_90_), 
	.A(prev_key1_reg[90]));
   DLY4X1 FE_PHC923_n1071 (.Y(FE_PHN923_n1071), 
	.A(FE_PHN4136_n1071));
   DLY4X1 FE_PHC922_prev_key1_reg_89_ (.Y(FE_PHN922_prev_key1_reg_89_), 
	.A(prev_key1_reg[89]));
   DLY4X1 FE_PHC921_prev_key1_reg_91_ (.Y(FE_PHN921_prev_key1_reg_91_), 
	.A(prev_key1_reg[91]));
   DLY4X1 FE_PHC919_prev_key1_reg_92_ (.Y(FE_PHN919_prev_key1_reg_92_), 
	.A(prev_key1_reg[92]));
   DLY4X1 FE_PHC917_key_mem_676_ (.Y(FE_PHN917_key_mem_676_), 
	.A(key_mem[676]));
   DLY4X1 FE_PHC916_n1600 (.Y(FE_PHN916_n1600), 
	.A(FE_PHN4012_n1600));
   DLY4X1 FE_PHC915_key_mem_371_ (.Y(FE_PHN915_key_mem_371_), 
	.A(key_mem[371]));
   DLY4X1 FE_PHC914_key_mem_652_ (.Y(FE_PHN914_key_mem_652_), 
	.A(key_mem[652]));
   DLY4X1 FE_PHC913_n2157 (.Y(FE_PHN913_n2157), 
	.A(FE_PHN4358_n2157));
   DLY4X1 FE_PHC912_rcon_reg_7_ (.Y(FE_PHN912_rcon_reg_7_), 
	.A(rcon_reg[7]));
   DLY4X1 FE_PHC896_prev_key1_reg_61_ (.Y(FE_PHN896_prev_key1_reg_61_), 
	.A(prev_key1_reg[61]));
   DLY4X1 FE_PHC827_n2122 (.Y(FE_PHN827_n2122), 
	.A(FE_PHN4051_n2122));
   DLY4X1 FE_PHC819_key_mem_1176_ (.Y(FE_PHN819_key_mem_1176_), 
	.A(key_mem[1176]));
   DLY4X1 FE_PHC817_key_mem_1240_ (.Y(FE_PHN817_key_mem_1240_), 
	.A(key_mem[1240]));
   DLY4X1 FE_PHC812_n1206 (.Y(FE_PHN812_n1206), 
	.A(FE_PHN4796_n1206));
   DLY4X1 FE_PHC811_key_mem_1247_ (.Y(FE_PHN811_key_mem_1247_), 
	.A(key_mem[1247]));
   DLY4X1 FE_PHC810_n1059 (.Y(FE_PHN810_n1059), 
	.A(FE_PHN4762_n1059));
   DLY4X1 FE_PHC808_key_mem_1182_ (.Y(FE_PHN808_key_mem_1182_), 
	.A(key_mem[1182]));
   DLY4X1 FE_PHC807_n1146 (.Y(FE_PHN807_n1146), 
	.A(FE_PHN4545_n1146));
   DLY4X1 FE_PHC806_n1317 (.Y(FE_PHN806_n1317), 
	.A(FE_PHN4670_n1317));
   DLY4X1 FE_PHC803_n1190 (.Y(FE_PHN803_n1190), 
	.A(FE_PHN4559_n1190));
   DLY4X1 FE_PHC802_key_mem_1273_ (.Y(FE_PHN802_key_mem_1273_), 
	.A(key_mem[1273]));
   DLY4X1 FE_PHC800_key_mem_1214_ (.Y(FE_PHN800_key_mem_1214_), 
	.A(key_mem[1214]));
   DLY4X1 FE_PHC798_key_mem_1166_ (.Y(FE_PHN798_key_mem_1166_), 
	.A(key_mem[1166]));
   DLY4X1 FE_PHC797_key_mem_1212_ (.Y(FE_PHN797_key_mem_1212_), 
	.A(key_mem[1212]));
   DLY4X1 FE_PHC796_n1342 (.Y(FE_PHN796_n1342), 
	.A(FE_PHN4343_n1342));
   DLY4X1 FE_PHC794_key_mem_1246_ (.Y(FE_PHN794_key_mem_1246_), 
	.A(key_mem[1246]));
   DLY4X1 FE_PHC792_key_mem_1277_ (.Y(FE_PHN792_key_mem_1277_), 
	.A(key_mem[1277]));
   DLY4X1 FE_PHC791_key_mem_1177_ (.Y(FE_PHN791_key_mem_1177_), 
	.A(key_mem[1177]));
   DLY4X1 FE_PHC789_n1205 (.Y(FE_PHN789_n1205), 
	.A(FE_PHN4707_n1205));
   DLY4X1 FE_PHC788_key_mem_1372_ (.Y(FE_PHN788_key_mem_1372_), 
	.A(key_mem[1372]));
   DLY4X1 FE_PHC786_key_mem_1208_ (.Y(FE_PHN786_key_mem_1208_), 
	.A(key_mem[1208]));
   DLY4X1 FE_PHC785_key_mem_1218_ (.Y(FE_PHN785_key_mem_1218_), 
	.A(key_mem[1218]));
   DLY4X1 FE_PHC783_key_mem_1209_ (.Y(FE_PHN783_key_mem_1209_), 
	.A(key_mem[1209]));
   DLY4X1 FE_PHC782_key_mem_1213_ (.Y(FE_PHN782_key_mem_1213_), 
	.A(key_mem[1213]));
   DLY4X1 FE_PHC780_key_mem_1276_ (.Y(FE_PHN780_key_mem_1276_), 
	.A(key_mem[1276]));
   DLY4X1 FE_PHC779_key_mem_1249_ (.Y(FE_PHN779_key_mem_1249_), 
	.A(key_mem[1249]));
   DLY4X1 FE_PHC777_key_mem_1234_ (.Y(FE_PHN777_key_mem_1234_), 
	.A(key_mem[1234]));
   DLY4X1 FE_PHC776_key_mem_1239_ (.Y(FE_PHN776_key_mem_1239_), 
	.A(key_mem[1239]));
   DLY4X1 FE_PHC775_key_mem_1156_ (.Y(FE_PHN775_key_mem_1156_), 
	.A(key_mem[1156]));
   DLY4X1 FE_PHC774_key_mem_1345_ (.Y(FE_PHN774_key_mem_1345_), 
	.A(key_mem[1345]));
   DLY4X1 FE_PHC773_key_mem_1245_ (.Y(FE_PHN773_key_mem_1245_), 
	.A(key_mem[1245]));
   DLY4X1 FE_PHC772_key_mem_760_ (.Y(FE_PHN772_key_mem_760_), 
	.A(key_mem[760]));
   DLY4X1 FE_PHC771_key_mem_1243_ (.Y(FE_PHN771_key_mem_1243_), 
	.A(key_mem[1243]));
   DLY4X1 FE_PHC770_key_mem_1241_ (.Y(FE_PHN770_key_mem_1241_), 
	.A(key_mem[1241]));
   DLY4X1 FE_PHC769_n1323 (.Y(FE_PHN769_n1323), 
	.A(n1323));
   DLY4X1 FE_PHC768_key_mem_1173_ (.Y(FE_PHN768_key_mem_1173_), 
	.A(key_mem[1173]));
   DLY4X1 FE_PHC767_key_mem_1242_ (.Y(FE_PHN767_key_mem_1242_), 
	.A(key_mem[1242]));
   DLY4X1 FE_PHC766_key_mem_1274_ (.Y(FE_PHN766_key_mem_1274_), 
	.A(key_mem[1274]));
   DLY4X1 FE_PHC765_key_mem_1211_ (.Y(FE_PHN765_key_mem_1211_), 
	.A(key_mem[1211]));
   DLY4X1 FE_PHC764_key_mem_287_ (.Y(FE_PHN764_key_mem_287_), 
	.A(key_mem[287]));
   DLY4X1 FE_PHC763_key_mem_275_ (.Y(FE_PHN763_key_mem_275_), 
	.A(key_mem[275]));
   DLY4X1 FE_PHC762_key_mem_767_ (.Y(FE_PHN762_key_mem_767_), 
	.A(key_mem[767]));
   DLY4X1 FE_PHC760_key_mem_1179_ (.Y(FE_PHN760_key_mem_1179_), 
	.A(key_mem[1179]));
   DLY4X1 FE_PHC758_key_mem_703_ (.Y(FE_PHN758_key_mem_703_), 
	.A(key_mem[703]));
   DLY4X1 FE_PHC757_prev_key1_reg_93_ (.Y(FE_PHN757_prev_key1_reg_93_), 
	.A(prev_key1_reg[93]));
   DLY4X1 FE_PHC756_key_mem_766_ (.Y(FE_PHN756_key_mem_766_), 
	.A(key_mem[766]));
   DLY4X1 FE_PHC755_key_mem_379_ (.Y(FE_PHN755_key_mem_379_), 
	.A(key_mem[379]));
   DLY4X1 FE_PHC754_key_mem_657_ (.Y(FE_PHN754_key_mem_657_), 
	.A(key_mem[657]));
   DLY4X1 FE_PHC748_keymem_sboxw_6_ (.Y(sboxw[6]), 
	.A(FE_PHN748_keymem_sboxw_6_));
   DLY4X1 FE_PHC747_n2364 (.Y(FE_PHN747_n2364), 
	.A(FE_PHN5006_n2364));
   DLY4X1 FE_PHC746_prev_key1_reg_58_ (.Y(FE_PHN746_prev_key1_reg_58_), 
	.A(prev_key1_reg[58]));
   DLY4X1 FE_PHC745_prev_key1_reg_59_ (.Y(FE_PHN745_prev_key1_reg_59_), 
	.A(prev_key1_reg[59]));
   DLY4X1 FE_PHC744_prev_key1_reg_57_ (.Y(FE_PHN744_prev_key1_reg_57_), 
	.A(prev_key1_reg[57]));
   DLY4X1 FE_PHC743_prev_key1_reg_63_ (.Y(FE_PHN743_prev_key1_reg_63_), 
	.A(prev_key1_reg[63]));
   DLY4X1 FE_PHC741_prev_key1_reg_60_ (.Y(FE_PHN741_prev_key1_reg_60_), 
	.A(prev_key1_reg[60]));
   DLY4X1 FE_PHC740_prev_key1_reg_62_ (.Y(FE_PHN740_prev_key1_reg_62_), 
	.A(prev_key1_reg[62]));
   DLY4X1 FE_PHC739_n1244 (.Y(FE_PHN739_n1244), 
	.A(FE_PHN4878_n1244));
   DLY4X1 FE_PHC738_n1365 (.Y(FE_PHN738_n1365), 
	.A(FE_PHN4724_n1365));
   DLY4X1 FE_PHC737_n1354 (.Y(FE_PHN737_n1354), 
	.A(FE_PHN4739_n1354));
   DLY4X1 FE_PHC736_n1219 (.Y(FE_PHN736_n1219), 
	.A(FE_PHN4637_n1219));
   DLY4X1 FE_PHC735_n1225 (.Y(FE_PHN735_n1225), 
	.A(FE_PHN4310_n1225));
   DLY4X1 FE_PHC734_n1345 (.Y(FE_PHN734_n1345), 
	.A(FE_PHN4519_n1345));
   DLY4X1 FE_PHC733_n1360 (.Y(FE_PHN733_n1360), 
	.A(FE_PHN4552_n1360));
   DLY4X1 FE_PHC732_n1343 (.Y(FE_PHN732_n1343), 
	.A(FE_PHN4429_n1343));
   DLY4X1 FE_PHC731_n953 (.Y(FE_PHN731_n953), 
	.A(FE_PHN4696_n953));
   DLY4X1 FE_PHC730_n1112 (.Y(FE_PHN730_n1112), 
	.A(FE_PHN4239_n1112));
   DLY4X1 FE_PHC728_n1236 (.Y(FE_PHN728_n1236), 
	.A(FE_PHN4240_n1236));
   DLY4X1 FE_PHC727_n968 (.Y(FE_PHN727_n968), 
	.A(FE_PHN4074_n968));
   DLY4X1 FE_PHC726_n1095 (.Y(FE_PHN726_n1095), 
	.A(FE_PHN4102_n1095));
   DLY4X1 FE_PHC724_n1107 (.Y(FE_PHN724_n1107), 
	.A(FE_PHN4262_n1107));
   DLY4X1 FE_PHC723_n1366 (.Y(FE_PHN723_n1366), 
	.A(FE_PHN4351_n1366));
   DLY4X1 FE_PHC722_n1335 (.Y(FE_PHN722_n1335), 
	.A(FE_PHN4151_n1335));
   DLY4X1 FE_PHC721_n1111 (.Y(FE_PHN721_n1111), 
	.A(FE_PHN4216_n1111));
   DLY4X1 FE_PHC720_n1088 (.Y(FE_PHN720_n1088), 
	.A(FE_PHN4129_n1088));
   DLY4X1 FE_PHC719_n978 (.Y(FE_PHN719_n978), 
	.A(FE_PHN4316_n978));
   DLY4X1 FE_PHC718_n962 (.Y(FE_PHN718_n962), 
	.A(FE_PHN3869_n962));
   DLY4X1 FE_PHC717_n987 (.Y(FE_PHN717_n987), 
	.A(n987));
   DLY4X1 FE_PHC716_n1105 (.Y(FE_PHN716_n1105), 
	.A(FE_PHN4350_n1105));
   DLY4X1 FE_PHC715_n2372 (.Y(FE_PHN715_n2372), 
	.A(FE_PHN3819_n2372));
   DLY4X1 FE_PHC714_n2374 (.Y(FE_PHN714_n2374), 
	.A(FE_PHN3858_n2374));
   DLY4X1 FE_PHC713_n1114 (.Y(FE_PHN713_n1114), 
	.A(FE_PHN3967_n1114));
   DLY4X1 FE_PHC712_n955 (.Y(FE_PHN712_n955), 
	.A(FE_PHN3956_n955));
   DLY4X1 FE_PHC710_n1364 (.Y(FE_PHN710_n1364), 
	.A(FE_PHN3782_n1364));
   DLY4X1 FE_PHC709_n985 (.Y(FE_PHN709_n985), 
	.A(FE_PHN3941_n985));
   DLY4X1 FE_PHC708_n975 (.Y(FE_PHN708_n975), 
	.A(FE_PHN4336_n975));
   DLY4X1 FE_PHC707_n1336 (.Y(FE_PHN707_n1336), 
	.A(FE_PHN4079_n1336));
   DLY4X1 FE_PHC706_n1102 (.Y(FE_PHN706_n1102), 
	.A(FE_PHN4253_n1102));
   DLY4X1 FE_PHC705_n629 (.Y(FE_PHN705_n629), 
	.A(n629));
   DLY4X1 FE_PHC700_key_mem_1265_ (.Y(FE_PHN700_key_mem_1265_), 
	.A(key_mem[1265]));
   DLY4X1 FE_PHC699_key_mem_1254_ (.Y(FE_PHN699_key_mem_1254_), 
	.A(key_mem[1254]));
   DLY4X1 FE_PHC698_key_mem_1172_ (.Y(FE_PHN698_key_mem_1172_), 
	.A(key_mem[1172]));
   DLY4X1 FE_PHC696_key_mem_1194_ (.Y(FE_PHN696_key_mem_1194_), 
	.A(key_mem[1194]));
   DLY4X1 FE_PHC694_key_mem_1232_ (.Y(FE_PHN694_key_mem_1232_), 
	.A(key_mem[1232]));
   DLY4X1 FE_PHC692_key_mem_1226_ (.Y(FE_PHN692_key_mem_1226_), 
	.A(key_mem[1226]));
   DLY4X1 FE_PHC691_key_mem_1248_ (.Y(FE_PHN691_key_mem_1248_), 
	.A(key_mem[1248]));
   DLY4X1 FE_PHC689_key_mem_1223_ (.Y(FE_PHN689_key_mem_1223_), 
	.A(key_mem[1223]));
   DLY4X1 FE_PHC688_key_mem_1252_ (.Y(FE_PHN688_key_mem_1252_), 
	.A(key_mem[1252]));
   DLY4X1 FE_PHC686_key_mem_1250_ (.Y(FE_PHN686_key_mem_1250_), 
	.A(key_mem[1250]));
   DLY4X1 FE_PHC684_key_mem_640_ (.Y(FE_PHN684_key_mem_640_), 
	.A(key_mem[640]));
   DLY4X1 FE_PHC683_key_mem_641_ (.Y(FE_PHN683_key_mem_641_), 
	.A(key_mem[641]));
   DLY4X1 FE_PHC646_n1308 (.Y(FE_PHN646_n1308), 
	.A(FE_PHN4936_n1308));
   DLY4X1 FE_PHC638_n1048 (.Y(FE_PHN638_n1048), 
	.A(FE_PHN4913_n1048));
   DLY4X1 FE_PHC635_n1373 (.Y(FE_PHN635_n1373), 
	.A(FE_PHN4433_n1373));
   DLY4X1 FE_PHC633_n1305 (.Y(FE_PHN633_n1305), 
	.A(FE_PHN4315_n1305));
   DLY4X1 FE_PHC632_n1175 (.Y(FE_PHN632_n1175), 
	.A(FE_PHN3992_n1175));
   DLY4X1 FE_PHC631_n917 (.Y(FE_PHN631_n917), 
	.A(n917));
   DLY4X1 FE_PHC628_n923 (.Y(FE_PHN628_n923), 
	.A(FE_PHN3884_n923));
   DLY4X1 FE_PHC627_n1768 (.Y(FE_PHN627_n1768), 
	.A(FE_PHN3885_n1768));
   DLY4X1 FE_PHC626_n1439 (.Y(FE_PHN626_n1439), 
	.A(FE_PHN3716_n1439));
   DLY4X1 FE_PHC625_n649 (.Y(FE_PHN625_n649), 
	.A(n649));
   DLY4X1 FE_PHC624_n551 (.Y(FE_PHN624_n551), 
	.A(n551));
   DLY4X1 FE_PHC623_n544 (.Y(FE_PHN623_n544), 
	.A(n544));
   DLY4X1 FE_PHC622_n543 (.Y(FE_PHN622_n543), 
	.A(n543));
   DLY4X1 FE_PHC621_n561 (.Y(FE_PHN621_n561), 
	.A(n561));
   DLY4X1 FE_PHC620_n554 (.Y(FE_PHN620_n554), 
	.A(n554));
   DLY4X1 FE_PHC619_n555 (.Y(FE_PHN619_n555), 
	.A(n555));
   DLY4X1 FE_PHC618_n562 (.Y(FE_PHN618_n562), 
	.A(n562));
   DLY4X1 FE_PHC617_n570 (.Y(FE_PHN617_n570), 
	.A(n570));
   DLY4X1 FE_PHC616_n553 (.Y(FE_PHN616_n553), 
	.A(n553));
   DLY4X1 FE_PHC615_n563 (.Y(FE_PHN615_n563), 
	.A(n563));
   DLY4X1 FE_PHC614_n556 (.Y(FE_PHN614_n556), 
	.A(n556));
   DLY4X1 FE_PHC613_n569 (.Y(FE_PHN613_n569), 
	.A(n569));
   DLY4X1 FE_PHC612_n572 (.Y(FE_PHN612_n572), 
	.A(n572));
   DLY4X1 FE_PHC611_n567 (.Y(FE_PHN611_n567), 
	.A(n567));
   DLY4X1 FE_PHC610_n573 (.Y(FE_PHN610_n573), 
	.A(n573));
   DLY4X1 FE_PHC609_n574 (.Y(FE_PHN609_n574), 
	.A(n574));
   DLY4X1 FE_PHC608_n564 (.Y(FE_PHN608_n564), 
	.A(n564));
   DLY4X1 FE_PHC607_n566 (.Y(FE_PHN607_n566), 
	.A(n566));
   DLY4X1 FE_PHC606_n571 (.Y(FE_PHN606_n571), 
	.A(n571));
   DLY4X1 FE_PHC605_n568 (.Y(FE_PHN605_n568), 
	.A(n568));
   DLY4X1 FE_PHC594_key_mem_1225_ (.Y(FE_PHN594_key_mem_1225_), 
	.A(key_mem[1225]));
   DLY4X1 FE_PHC593_n1381 (.Y(FE_PHN593_n1381), 
	.A(FE_PHN4606_n1381));
   DLY4X1 FE_PHC592_key_mem_1390_ (.Y(FE_PHN592_key_mem_1390_), 
	.A(key_mem[1390]));
   DLY4X1 FE_PHC591_key_mem_1230_ (.Y(FE_PHN591_key_mem_1230_), 
	.A(key_mem[1230]));
   DLY4X1 FE_PHC590_n1389 (.Y(FE_PHN590_n1389), 
	.A(FE_PHN4306_n1389));
   DLY4X1 FE_PHC589_n1082 (.Y(FE_PHN589_n1082), 
	.A(FE_PHN4295_n1082));
   DLY4X1 FE_PHC588_n1259 (.Y(FE_PHN588_n1259), 
	.A(n1259));
   DLY4X1 FE_PHC587_key_mem_1161_ (.Y(FE_PHN587_key_mem_1161_), 
	.A(key_mem[1161]));
   DLY4X1 FE_PHC586_n1132 (.Y(FE_PHN586_n1132), 
	.A(FE_PHN4569_n1132));
   DLY4X1 FE_PHC585_key_mem_1175_ (.Y(FE_PHN585_key_mem_1175_), 
	.A(key_mem[1175]));
   DLY4X1 FE_PHC584_key_mem_1159_ (.Y(FE_PHN584_key_mem_1159_), 
	.A(key_mem[1159]));
   DLY4X1 FE_PHC583_key_mem_1257_ (.Y(FE_PHN583_key_mem_1257_), 
	.A(key_mem[1257]));
   DLY4X1 FE_PHC582_key_mem_1170_ (.Y(FE_PHN582_key_mem_1170_), 
	.A(key_mem[1170]));
   DLY4X1 FE_PHC581_n1004 (.Y(FE_PHN581_n1004), 
	.A(FE_PHN4544_n1004));
   DLY4X1 FE_PHC580_key_mem_743_ (.Y(FE_PHN580_key_mem_743_), 
	.A(key_mem[743]));
   DLY3X1 FE_PHC579_n650 (.Y(FE_PHN579_n650), 
	.A(n650));
   DLY4X1 FE_PHC578_n600 (.Y(FE_PHN578_n600), 
	.A(n600));
   DLY4X1 FE_PHC577_n593 (.Y(FE_PHN577_n593), 
	.A(n593));
   DLY4X1 FE_PHC576_n584 (.Y(FE_PHN576_n584), 
	.A(n584));
   DLY4X1 FE_PHC575_n594 (.Y(FE_PHN575_n594), 
	.A(n594));
   DLY4X1 FE_PHC574_n583 (.Y(FE_PHN574_n583), 
	.A(n583));
   DLY4X1 FE_PHC573_n654 (.Y(FE_PHN573_n654), 
	.A(n654));
   DLY4X1 FE_PHC572_n664 (.Y(FE_PHN572_n664), 
	.A(n664));
   DLY4X1 FE_PHC571_n656 (.Y(FE_PHN571_n656), 
	.A(n656));
   DLY4X1 FE_PHC570_n653 (.Y(FE_PHN570_n653), 
	.A(n653));
   DLY4X1 FE_PHC569_n651 (.Y(FE_PHN569_n651), 
	.A(n651));
   DLY4X1 FE_PHC568_n550 (.Y(FE_PHN568_n550), 
	.A(n550));
   DLY4X1 FE_PHC567_n549 (.Y(FE_PHN567_n549), 
	.A(n549));
   DLY4X1 FE_PHC566_n665 (.Y(FE_PHN566_n665), 
	.A(n665));
   DLY4X1 FE_PHC565_n596 (.Y(FE_PHN565_n596), 
	.A(n596));
   DLY4X1 FE_PHC564_n648 (.Y(FE_PHN564_n648), 
	.A(n648));
   DLY4X1 FE_PHC563_n667 (.Y(FE_PHN563_n667), 
	.A(n667));
   DLY4X1 FE_PHC562_n666 (.Y(FE_PHN562_n666), 
	.A(n666));
   DLY4X1 FE_PHC561_n601 (.Y(FE_PHN561_n601), 
	.A(n601));
   DLY4X1 FE_PHC560_n658 (.Y(FE_PHN560_n658), 
	.A(n658));
   DLY4X1 FE_PHC559_n598 (.Y(FE_PHN559_n598), 
	.A(n598));
   DLY4X1 FE_PHC558_n652 (.Y(FE_PHN558_n652), 
	.A(n652));
   DLY4X1 FE_PHC557_n602 (.Y(FE_PHN557_n602), 
	.A(n602));
   DLY4X1 FE_PHC556_n595 (.Y(FE_PHN556_n595), 
	.A(n595));
   DLY4X1 FE_PHC555_n605 (.Y(FE_PHN555_n605), 
	.A(n605));
   DLY4X1 FE_PHC554_n659 (.Y(FE_PHN554_n659), 
	.A(n659));
   DLY4X1 FE_PHC553_n670 (.Y(FE_PHN553_n670), 
	.A(n670));
   DLY4X1 FE_PHC552_n657 (.Y(FE_PHN552_n657), 
	.A(n657));
   DLY4X1 FE_PHC551_n545 (.Y(FE_PHN551_n545), 
	.A(n545));
   DLY4X1 FE_PHC550_n668 (.Y(FE_PHN550_n668), 
	.A(n668));
   DLY4X1 FE_PHC549_n587 (.Y(FE_PHN549_n587), 
	.A(n587));
   DLY4X1 FE_PHC548_n546 (.Y(FE_PHN548_n546), 
	.A(n546));
   DLY4X1 FE_PHC547_n580 (.Y(FE_PHN547_n580), 
	.A(n580));
   DLY4X1 FE_PHC546_n603 (.Y(FE_PHN546_n603), 
	.A(n603));
   DLY4X1 FE_PHC545_n599 (.Y(FE_PHN545_n599), 
	.A(n599));
   DLY4X1 FE_PHC544_n547 (.Y(FE_PHN544_n547), 
	.A(n547));
   DLY4X1 FE_PHC543_n588 (.Y(FE_PHN543_n588), 
	.A(n588));
   DLY4X1 FE_PHC542_n586 (.Y(FE_PHN542_n586), 
	.A(n586));
   DLY4X1 FE_PHC541_n660 (.Y(FE_PHN541_n660), 
	.A(n660));
   DLY4X1 FE_PHC540_n606 (.Y(FE_PHN540_n606), 
	.A(n606));
   DLY4X1 FE_PHC539_n585 (.Y(FE_PHN539_n585), 
	.A(n585));
   DLY4X1 FE_PHC538_n604 (.Y(FE_PHN538_n604), 
	.A(n604));
   DLY4X1 FE_PHC537_n669 (.Y(FE_PHN537_n669), 
	.A(n669));
   DLY4X1 FE_PHC432_key_mem_1256_ (.Y(FE_PHN432_key_mem_1256_), 
	.A(key_mem[1256]));
   DLY4X1 FE_PHC431_key_mem_1224_ (.Y(FE_PHN431_key_mem_1224_), 
	.A(key_mem[1224]));
   DLY4X1 FE_PHC430_key_mem_1167_ (.Y(FE_PHN430_key_mem_1167_), 
	.A(key_mem[1167]));
   DLY4X1 FE_PHC429_key_mem_1162_ (.Y(FE_PHN429_key_mem_1162_), 
	.A(key_mem[1162]));
   DLY4X1 FE_PHC428_n1161 (.Y(FE_PHN428_n1161), 
	.A(FE_PHN4170_n1161));
   DLY4X1 FE_PHC427_key_mem_1258_ (.Y(FE_PHN427_key_mem_1258_), 
	.A(key_mem[1258]));
   DLY4X1 FE_PHC426_key_mem_1184_ (.Y(FE_PHN426_key_mem_1184_), 
	.A(key_mem[1184]));
   DLY4X1 FE_PHC425_key_mem_1264_ (.Y(FE_PHN425_key_mem_1264_), 
	.A(key_mem[1264]));
   DLY4X1 FE_PHC424_key_mem_367_ (.Y(FE_PHN424_key_mem_367_), 
	.A(key_mem[367]));
   DLY4X1 FE_PHC423_n607 (.Y(FE_PHN423_n607), 
	.A(n607));
   DLY4X1 FE_PHC422_n608 (.Y(FE_PHN422_n608), 
	.A(n608));
   DLY4X1 FE_PHC421_n590 (.Y(FE_PHN421_n590), 
	.A(n590));
   DLY4X1 FE_PHC420_n592 (.Y(FE_PHN420_n592), 
	.A(n592));
   DLY4X1 FE_PHC419_n589 (.Y(FE_PHN419_n589), 
	.A(n589));
   DLY4X1 FE_PHC418_n548 (.Y(FE_PHN418_n548), 
	.A(n548));
   DLY4X1 FE_PHC417_n591 (.Y(FE_PHN417_n591), 
	.A(n591));
   DLY4X1 FE_PHC416_n597 (.Y(FE_PHN416_n597), 
	.A(n597));
   DLY4X1 FE_PHC411_n6 (.Y(FE_PHN411_n6), 
	.A(n6));
   DLY4X1 FE_PHC409_n624 (.Y(FE_PHN409_n624), 
	.A(n624));
   DLY4X1 FE_PHC408_n640 (.Y(FE_PHN408_n640), 
	.A(n640));
   DLY4X1 FE_PHC407_n645 (.Y(FE_PHN407_n645), 
	.A(n645));
   DLY4X1 FE_PHC406_n646 (.Y(FE_PHN406_n646), 
	.A(n646));
   DLY4X1 FE_PHC405_n613 (.Y(FE_PHN405_n613), 
	.A(n613));
   DLY4X1 FE_PHC404_n614 (.Y(FE_PHN404_n614), 
	.A(n614));
   DLY4X1 FE_PHC403_n622 (.Y(FE_PHN403_n622), 
	.A(n622));
   DLY4X1 FE_PHC402_n621 (.Y(FE_PHN402_n621), 
	.A(n621));
   DLY4X1 FE_PHC401_n639 (.Y(FE_PHN401_n639), 
	.A(n639));
   DLY4X1 FE_PHC400_n641 (.Y(FE_PHN400_n641), 
	.A(n641));
   DLY4X1 FE_PHC399_n643 (.Y(FE_PHN399_n643), 
	.A(n643));
   DLY4X1 FE_PHC398_n627 (.Y(FE_PHN398_n627), 
	.A(n627));
   DLY4X1 FE_PHC397_n642 (.Y(FE_PHN397_n642), 
	.A(n642));
   DLY4X1 FE_PHC396_n632 (.Y(FE_PHN396_n632), 
	.A(n632));
   DLY4X1 FE_PHC395_n644 (.Y(FE_PHN395_n644), 
	.A(n644));
   DLY4X1 FE_PHC394_n634 (.Y(FE_PHN394_n634), 
	.A(n634));
   DLY4X1 FE_PHC393_n609 (.Y(FE_PHN393_n609), 
	.A(n609));
   DLY4X1 FE_PHC392_n610 (.Y(FE_PHN392_n610), 
	.A(n610));
   DLY4X1 FE_PHC391_n633 (.Y(FE_PHN391_n633), 
	.A(n633));
   DLY4X1 FE_PHC390_n628 (.Y(FE_PHN390_n628), 
	.A(n628));
   DLY4X1 FE_PHC389_n618 (.Y(FE_PHN389_n618), 
	.A(n618));
   DLY4X1 FE_PHC388_n626 (.Y(FE_PHN388_n626), 
	.A(n626));
   DLY4X1 FE_PHC387_n625 (.Y(FE_PHN387_n625), 
	.A(n625));
   DLY4X1 FE_PHC386_n611 (.Y(FE_PHN386_n611), 
	.A(n611));
   DLY4X1 FE_PHC385_n617 (.Y(FE_PHN385_n617), 
	.A(n617));
   DLY4X1 FE_PHC384_n620 (.Y(FE_PHN384_n620), 
	.A(n620));
   DLY4X1 FE_PHC383_n638 (.Y(FE_PHN383_n638), 
	.A(n638));
   DLY4X1 FE_PHC382_n619 (.Y(FE_PHN382_n619), 
	.A(n619));
   DLY4X1 FE_PHC381_n636 (.Y(FE_PHN381_n636), 
	.A(n636));
   DLY4X1 FE_PHC380_n637 (.Y(FE_PHN380_n637), 
	.A(n637));
   DLY4X1 FE_PHC379_n635 (.Y(FE_PHN379_n635), 
	.A(n635));
   DLY4X1 FE_PHC360_prev_key1_reg_86_ (.Y(FE_PHN360_prev_key1_reg_86_), 
	.A(prev_key1_reg[86]));
   DLY4X1 FE_PHC359_prev_key1_reg_87_ (.Y(FE_PHN359_prev_key1_reg_87_), 
	.A(prev_key1_reg[87]));
   DLY4X1 FE_PHC357_key_mem_1154_ (.Y(FE_PHN357_key_mem_1154_), 
	.A(key_mem[1154]));
   DLY4X1 FE_PHC349_n581 (.Y(FE_PHN349_n581), 
	.A(n581));
   DLY4X1 FE_PHC348_n647 (.Y(FE_PHN348_n647), 
	.A(n647));
   DLY4X1 FE_PHC347_n582 (.Y(FE_PHN347_n582), 
	.A(n582));
   DLY4X1 FE_PHC346_n579 (.Y(FE_PHN346_n579), 
	.A(n579));
   DLY4X1 FE_PHC345_n578 (.Y(FE_PHN345_n578), 
	.A(n578));
   DLY4X1 FE_PHC344_n576 (.Y(FE_PHN344_n576), 
	.A(n576));
   DLY4X1 FE_PHC343_n577 (.Y(FE_PHN343_n577), 
	.A(n577));
   DLY4X1 FE_PHC342_n575 (.Y(FE_PHN342_n575), 
	.A(n575));
   DLY4X1 FE_PHC327_n655 (.Y(FE_PHN327_n655), 
	.A(n655));
   DLY4X1 FE_PHC326_n612 (.Y(FE_PHN326_n612), 
	.A(n612));
   DLY4X1 FE_PHC325_n662 (.Y(FE_PHN325_n662), 
	.A(n662));
   DLY4X1 FE_PHC324_n663 (.Y(FE_PHN324_n663), 
	.A(n663));
   DLY4X1 FE_PHC323_n661 (.Y(FE_PHN323_n661), 
	.A(n661));
   DLY4X1 FE_PHC290_key_mem_ctrl_reg_0_ (.Y(FE_PHN290_key_mem_ctrl_reg_0_), 
	.A(key_mem_ctrl_reg[0]));
   DLY4X1 FE_PHC283_n2433 (.Y(FE_PHN283_n2433), 
	.A(n2433));
   DLY4X1 FE_PHC265_keymem_sboxw_7_ (.Y(sboxw[7]), 
	.A(FE_PHN265_keymem_sboxw_7_));
   DLY4X1 FE_PHC254_n689 (.Y(FE_PHN254_n689), 
	.A(n689));
   DLY4X1 FE_PHC198_round_ctr_reg_0_ (.Y(FE_PHN198_round_ctr_reg_0_), 
	.A(round_ctr_reg[0]));
   DLY4X1 FE_PHC178_round_ctr_reg_2_ (.Y(FE_PHN178_round_ctr_reg_2_), 
	.A(round_ctr_reg[2]));
   DLY4X1 FE_PHC155_n3 (.Y(FE_PHN155_n3), 
	.A(n3));
   DLY4X1 FE_PHC120_key_mem_ctrl_reg_1_ (.Y(FE_PHN120_key_mem_ctrl_reg_1_), 
	.A(key_mem_ctrl_reg[1]));
   DLY4X1 FE_PHC116_round_ctr_reg_3_ (.Y(FE_PHN116_round_ctr_reg_3_), 
	.A(round_ctr_reg[3]));
   DLY4X1 FE_PHC112_round_ctr_reg_1_ (.Y(FE_PHN112_round_ctr_reg_1_), 
	.A(round_ctr_reg[1]));
   CLKBUFX4 FE_OFC109_n23 (.Y(FE_OFN109_n23), 
	.A(n23));
   CLKBUFX2 FE_OFC108_n21 (.Y(FE_OFN108_n21), 
	.A(n21));
   CLKBUFX2 FE_OFC107_n21 (.Y(FE_OFN107_n21), 
	.A(n21));
   CLKBUFX4 FE_OFC106_n22 (.Y(FE_OFN106_n22), 
	.A(n22));
   CLKBUFX4 FE_OFC105_n2763 (.Y(FE_OFN105_n2763), 
	.A(n2769));
   CLKBUFX4 FE_OFC104_n27 (.Y(FE_OFN104_n27), 
	.A(FE_OFN103_n27));
   CLKBUFX3 FE_OFC103_n27 (.Y(FE_OFN103_n27), 
	.A(n27));
   CLKBUFX4 FE_OFC102_n31 (.Y(FE_OFN102_n31), 
	.A(n31));
   CLKBUFX4 FE_OFC101_n30 (.Y(FE_OFN101_n30), 
	.A(n30));
   CLKBUFX3 FE_OFC100_n2800 (.Y(FE_OFN100_n2800), 
	.A(n2800));
   CLKBUFX4 FE_OFC99_n2811 (.Y(FE_OFN99_n2811), 
	.A(n2817));
   CLKBUFX2 FE_OFC96_n674 (.Y(FE_OFN96_n674), 
	.A(FE_OFN93_n674));
   CLKINVX3 FE_OFC95_n674 (.Y(FE_OFN95_n674), 
	.A(FE_OFN92_n674));
   CLKINVX2 FE_OFC94_n674 (.Y(FE_OFN94_n674), 
	.A(FE_OFN92_n674));
   CLKINVX2 FE_OFC93_n674 (.Y(FE_OFN93_n674), 
	.A(FE_OFN92_n674));
   INVX1 FE_OFC92_n674 (.Y(FE_OFN92_n674), 
	.A(n674));
   CLKBUFX3 FE_OFC91_n690 (.Y(FE_OFN91_n690), 
	.A(FE_OFN90_n690));
   CLKBUFX3 FE_OFC90_n690 (.Y(FE_OFN90_n690), 
	.A(n690));
   CLKBUFX2 FE_OFC89_n1 (.Y(FE_OFN89_n1), 
	.A(FE_OFN87_n1));
   CLKBUFX2 FE_OFC88_n1 (.Y(FE_OFN88_n1), 
	.A(FE_OFN86_n1));
   CLKINVX2 FE_OFC87_n1 (.Y(FE_OFN87_n1), 
	.A(FE_OFN84_n1));
   CLKINVX3 FE_OFC86_n1 (.Y(FE_OFN86_n1), 
	.A(FE_OFN84_n1));
   INVX2 FE_OFC85_n1 (.Y(FE_OFN85_n1), 
	.A(FE_OFN84_n1));
   INVX1 FE_OFC84_n1 (.Y(FE_OFN84_n1), 
	.A(n1));
   CLKINVX2 FE_OFC83_n672 (.Y(FE_OFN83_n672), 
	.A(FE_OFN79_n672));
   CLKINVX3 FE_OFC82_n672 (.Y(FE_OFN82_n672), 
	.A(FE_OFN79_n672));
   INVX2 FE_OFC81_n672 (.Y(FE_OFN81_n672), 
	.A(FE_OFN79_n672));
   CLKINVX2 FE_OFC80_n672 (.Y(FE_OFN80_n672), 
	.A(FE_OFN79_n672));
   INVX1 FE_OFC79_n672 (.Y(FE_OFN79_n672), 
	.A(n672));
   CLKBUFX3 FE_OFC78_n676 (.Y(FE_OFN78_n676), 
	.A(FE_OFN77_n676));
   CLKBUFX3 FE_OFC77_n676 (.Y(FE_OFN77_n676), 
	.A(n676));
   CLKBUFX2 FE_OFC76_n676 (.Y(FE_OFN76_n676), 
	.A(n676));
   CLKINVX3 FE_OFC57_reset_n (.Y(FE_OFN57_reset_n), 
	.A(FE_OFN48_reset_n));
   CLKINVX3 FE_OFC41_reset_n (.Y(FE_OFN41_reset_n), 
	.A(reset_n));
   INVX1 FE_OFC36_reset_n (.Y(FE_OFN36_reset_n), 
	.A(reset_n));
   CLKBUFX2 FE_OFC33_n683 (.Y(FE_OFN33_n683), 
	.A(FE_OFN32_n683));
   CLKBUFX2 FE_OFC32_n683 (.Y(FE_OFN32_n683), 
	.A(FE_OFN31_n683));
   CLKBUFX2 FE_OFC31_n683 (.Y(FE_OFN31_n683), 
	.A(n683));
   CLKBUFX2 FE_OFC30_n687 (.Y(FE_OFN30_n687), 
	.A(FE_OFN29_n687));
   CLKBUFX2 FE_OFC29_n687 (.Y(FE_OFN29_n687), 
	.A(n687));
   CLKBUFX2 FE_OFC28_n687 (.Y(FE_OFN28_n687), 
	.A(n687));
   CLKBUFX3 FE_OFC27_n685 (.Y(FE_OFN27_n685), 
	.A(FE_OFN25_n685));
   CLKBUFX2 FE_OFC26_n685 (.Y(FE_OFN26_n685), 
	.A(n685));
   CLKBUFX2 FE_OFC25_n685 (.Y(FE_OFN25_n685), 
	.A(n685));
   BUFX1 FE_OFC24_n685 (.Y(FE_OFN24_n685), 
	.A(n685));
   CLKINVX2 FE_OFC23_n681 (.Y(FE_OFN23_n681), 
	.A(FE_OFN19_n681));
   CLKINVX2 FE_OFC22_n681 (.Y(FE_OFN22_n681), 
	.A(FE_OFN19_n681));
   INVX1 FE_OFC21_n681 (.Y(FE_OFN21_n681), 
	.A(FE_OFN19_n681));
   CLKINVX2 FE_OFC20_n681 (.Y(FE_OFN20_n681), 
	.A(FE_OFN19_n681));
   INVX1 FE_OFC19_n681 (.Y(FE_OFN19_n681), 
	.A(n681));
   CLKBUFX2 FE_OFC18_n678 (.Y(FE_OFN18_n678), 
	.A(FE_OFN15_n678));
   CLKBUFX2 FE_OFC17_n678 (.Y(FE_OFN17_n678), 
	.A(FE_OFN15_n678));
   CLKBUFX2 FE_OFC16_n678 (.Y(FE_OFN16_n678), 
	.A(FE_OFN15_n678));
   CLKBUFX3 FE_OFC15_n678 (.Y(FE_OFN15_n678), 
	.A(n678));
   CLKINVX2 FE_OFC14_n688 (.Y(FE_OFN14_n688), 
	.A(FE_OFN10_n688));
   CLKINVX2 FE_OFC13_n688 (.Y(FE_OFN13_n688), 
	.A(FE_OFN10_n688));
   INVX1 FE_OFC12_n688 (.Y(FE_OFN12_n688), 
	.A(FE_OFN10_n688));
   CLKINVX3 FE_OFC11_n688 (.Y(FE_OFN11_n688), 
	.A(FE_OFN10_n688));
   INVX1 FE_OFC10_n688 (.Y(FE_OFN10_n688), 
	.A(n688));
   CLKBUFX2 FE_OFC9_n684 (.Y(FE_OFN9_n684), 
	.A(FE_OFN7_n684));
   CLKBUFX2 FE_OFC8_n684 (.Y(FE_OFN8_n684), 
	.A(FE_OFN6_n684));
   CLKBUFX2 FE_OFC7_n684 (.Y(FE_OFN7_n684), 
	.A(FE_OFN6_n684));
   CLKBUFX2 FE_OFC6_n684 (.Y(FE_OFN6_n684), 
	.A(n684));
   CLKINVX2 FE_OFC5_n682 (.Y(FE_OFN5_n682), 
	.A(FE_OFN1_n682));
   CLKINVX2 FE_OFC4_n682 (.Y(FE_OFN4_n682), 
	.A(FE_OFN1_n682));
   INVX1 FE_OFC3_n682 (.Y(FE_OFN3_n682), 
	.A(FE_OFN1_n682));
   CLKINVX2 FE_OFC2_n682 (.Y(FE_OFN2_n682), 
	.A(FE_OFN1_n682));
   INVX1 FE_OFC1_n682 (.Y(FE_OFN1_n682), 
	.A(n682));
   NAND2X1 U1302 (.Y(n678), 
	.B(n680), 
	.A(n679));
   NAND4X1 U1431 (.Y(n681), 
	.D(n2874), 
	.C(FE_PHN198_round_ctr_reg_0_), 
	.B(FE_PHN178_round_ctr_reg_2_), 
	.A(n679));
   NAND3BX1 U1560 (.Y(n682), 
	.C(n680), 
	.B(FE_PHN112_round_ctr_reg_1_), 
	.AN(n683));
   OR3XL U1690 (.Y(n684), 
	.C(n2873), 
	.B(n683), 
	.A(n677));
   NAND2X2 U1819 (.Y(n685), 
	.B(FE_PHN411_n6), 
	.A(n686));
   NAND2X2 U1948 (.Y(n687), 
	.B(FE_PHN198_round_ctr_reg_0_), 
	.A(n686));
   OR2X2 U2079 (.Y(n688), 
	.B(n683), 
	.A(FE_PHN254_n689));
   NAND2X2 U2515 (.Y(n683), 
	.B(FE_OFN39_reset_n), 
	.A(FE_PHN155_n3));
   DFFHQX1 key_mem_reg_6__112_ (.Q(key_mem[624]), 
	.D(FE_PHN1759_n1668), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_6__111_ (.Q(key_mem[623]), 
	.D(FE_PHN2167_n1669), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_6__110_ (.Q(key_mem[622]), 
	.D(FE_PHN2496_n1670), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_6__109_ (.Q(key_mem[621]), 
	.D(FE_PHN1649_n1671), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_6__106_ (.Q(key_mem[618]), 
	.D(FE_PHN2350_n1674), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_6__104_ (.Q(key_mem[616]), 
	.D(FE_PHN2572_n1676), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_6__80_ (.Q(key_mem[592]), 
	.D(FE_PHN2420_n1683), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_6__79_ (.Q(key_mem[591]), 
	.D(FE_PHN2314_n1684), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_6__78_ (.Q(key_mem[590]), 
	.D(FE_PHN2246_n1685), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_6__77_ (.Q(key_mem[589]), 
	.D(FE_PHN2514_n1686), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_6__74_ (.Q(key_mem[586]), 
	.D(FE_PHN2559_n1689), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_6__72_ (.Q(key_mem[584]), 
	.D(FE_PHN2061_n1691), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_6__64_ (.Q(key_mem[576]), 
	.D(FE_PHN2523_n1699), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_6__48_ (.Q(key_mem[560]), 
	.D(FE_PHN2165_n1715), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_6__47_ (.Q(key_mem[559]), 
	.D(FE_PHN2575_n1716), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_6__46_ (.Q(key_mem[558]), 
	.D(FE_PHN2100_n1717), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_6__45_ (.Q(key_mem[557]), 
	.D(FE_PHN2122_n1718), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_6__42_ (.Q(key_mem[554]), 
	.D(FE_PHN2267_n1721), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_6__40_ (.Q(key_mem[552]), 
	.D(FE_PHN2437_n1723), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_6__32_ (.Q(key_mem[544]), 
	.D(FE_PHN2501_n1731), 
	.CK(clk));
   DFFHQX1 key_mem_reg_6__16_ (.Q(key_mem[528]), 
	.D(FE_PHN2473_n1747), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_6__15_ (.Q(key_mem[527]), 
	.D(FE_PHN2425_n1748), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_6__14_ (.Q(key_mem[526]), 
	.D(FE_PHN2635_n1749), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_6__13_ (.Q(key_mem[525]), 
	.D(FE_PHN1597_n1750), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_6__10_ (.Q(key_mem[522]), 
	.D(FE_PHN2068_n1753), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_6__8_ (.Q(key_mem[520]), 
	.D(FE_PHN2366_n1755), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_6__0_ (.Q(key_mem[512]), 
	.D(FE_PHN2055_n1763), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_6__96_ (.Q(key_mem[608]), 
	.D(FE_PHN1040_n1766), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_9__112_ (.Q(key_mem[240]), 
	.D(FE_PHN2341_n2052), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_9__111_ (.Q(key_mem[239]), 
	.D(FE_PHN2324_n2053), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_9__110_ (.Q(key_mem[238]), 
	.D(FE_PHN2188_n2054), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_9__109_ (.Q(key_mem[237]), 
	.D(FE_PHN2239_n2055), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_9__106_ (.Q(key_mem[234]), 
	.D(FE_PHN1612_n2058), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_9__104_ (.Q(key_mem[232]), 
	.D(FE_PHN2658_n2060), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_9__64_ (.Q(key_mem[192]), 
	.D(FE_PHN2361_n2071), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_9__48_ (.Q(key_mem[176]), 
	.D(FE_PHN2403_n2087), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_9__47_ (.Q(key_mem[175]), 
	.D(FE_PHN2057_n2088), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_9__46_ (.Q(key_mem[174]), 
	.D(FE_PHN2074_n2089), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_9__45_ (.Q(key_mem[173]), 
	.D(FE_PHN2245_n2090), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_9__42_ (.Q(key_mem[170]), 
	.D(FE_PHN2276_n2093), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_9__40_ (.Q(key_mem[168]), 
	.D(FE_PHN2293_n2095), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_9__32_ (.Q(key_mem[160]), 
	.D(FE_PHN2453_n2103), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_9__16_ (.Q(key_mem[144]), 
	.D(FE_PHN2667_n2119), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_9__15_ (.Q(key_mem[143]), 
	.D(FE_PHN2187_n2120), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_9__14_ (.Q(key_mem[142]), 
	.D(FE_PHN2138_n2121), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_9__13_ (.Q(key_mem[141]), 
	.D(FE_PHN827_n2122), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_9__10_ (.Q(key_mem[138]), 
	.D(FE_PHN1628_n2125), 
	.CK(clk_48Mhz__L6_N21));
   DFFHQX1 key_mem_reg_9__8_ (.Q(key_mem[136]), 
	.D(FE_PHN2355_n2127), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_9__0_ (.Q(key_mem[128]), 
	.D(FE_PHN2449_n2135), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_9__96_ (.Q(key_mem[224]), 
	.D(FE_PHN2071_n2138), 
	.CK(clk));
   DFFHQX1 key_mem_reg_9__80_ (.Q(key_mem[208]), 
	.D(FE_PHN2217_n2154), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_9__79_ (.Q(key_mem[207]), 
	.D(FE_PHN2287_n2155), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_9__78_ (.Q(key_mem[206]), 
	.D(FE_PHN2334_n2156), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_9__77_ (.Q(key_mem[205]), 
	.D(FE_PHN913_n2157), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_9__74_ (.Q(key_mem[202]), 
	.D(FE_PHN2144_n2160), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_9__72_ (.Q(key_mem[200]), 
	.D(FE_PHN2452_n2162), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_6__122_ (.Q(key_mem[634]), 
	.D(FE_PHN1467_n1658), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_9__122_ (.Q(key_mem[250]), 
	.D(FE_PHN1497_n2042), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_6__90_ (.Q(key_mem[602]), 
	.D(FE_PHN2450_n1772), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_9__90_ (.Q(key_mem[218]), 
	.D(FE_PHN1488_n2144), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_6__58_ (.Q(key_mem[570]), 
	.D(FE_PHN2172_n1705), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_9__58_ (.Q(key_mem[186]), 
	.D(FE_PHN1669_n2077), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_6__26_ (.Q(key_mem[538]), 
	.D(FE_PHN1474_n1737), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_9__26_ (.Q(key_mem[154]), 
	.D(FE_PHN2585_n2109), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_6__125_ (.Q(key_mem[637]), 
	.D(FE_PHN1675_n1655), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_9__125_ (.Q(key_mem[253]), 
	.D(FE_PHN2598_n2039), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_6__93_ (.Q(key_mem[605]), 
	.D(FE_PHN2043_n1769), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 key_mem_reg_9__93_ (.Q(key_mem[221]), 
	.D(FE_PHN2132_n2141), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 key_mem_reg_6__61_ (.Q(key_mem[573]), 
	.D(FE_PHN2422_n1702), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_9__61_ (.Q(key_mem[189]), 
	.D(FE_PHN2294_n2074), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_6__29_ (.Q(key_mem[541]), 
	.D(FE_PHN1708_n1734), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_9__29_ (.Q(key_mem[157]), 
	.D(FE_PHN1478_n2106), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_6__126_ (.Q(key_mem[638]), 
	.D(FE_PHN2396_n1654), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_9__126_ (.Q(key_mem[254]), 
	.D(FE_PHN2655_n2038), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_6__94_ (.Q(key_mem[606]), 
	.D(FE_PHN627_n1768), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 key_mem_reg_9__94_ (.Q(key_mem[222]), 
	.D(FE_PHN2261_n2140), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_6__62_ (.Q(key_mem[574]), 
	.D(FE_PHN2464_n1701), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_9__62_ (.Q(key_mem[190]), 
	.D(FE_PHN2045_n2073), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_6__30_ (.Q(key_mem[542]), 
	.D(FE_PHN2128_n1733), 
	.CK(clk_48Mhz__L6_N47));
   DFFHQX1 key_mem_reg_9__30_ (.Q(key_mem[158]), 
	.D(FE_PHN2076_n2105), 
	.CK(clk_48Mhz__L6_N47));
   DFFHQX1 key_mem_reg_6__120_ (.Q(key_mem[632]), 
	.D(FE_PHN1604_n1660), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_9__120_ (.Q(key_mem[248]), 
	.D(FE_PHN2053_n2044), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_6__88_ (.Q(key_mem[600]), 
	.D(FE_PHN2150_n1774), 
	.CK(clk_48Mhz__L6_N23));
   DFFHQX1 key_mem_reg_9__88_ (.Q(key_mem[216]), 
	.D(FE_PHN2113_n2146), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 key_mem_reg_6__56_ (.Q(key_mem[568]), 
	.D(FE_PHN2423_n1707), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_9__56_ (.Q(key_mem[184]), 
	.D(FE_PHN2084_n2079), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_6__24_ (.Q(key_mem[536]), 
	.D(FE_PHN1551_n1739), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_9__24_ (.Q(key_mem[152]), 
	.D(FE_PHN2649_n2111), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_6__127_ (.Q(key_mem[639]), 
	.D(FE_PHN2135_n1653), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_9__127_ (.Q(key_mem[255]), 
	.D(FE_PHN2477_n2037), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_6__95_ (.Q(key_mem[607]), 
	.D(FE_PHN2318_n1767), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_9__95_ (.Q(key_mem[223]), 
	.D(FE_PHN2534_n2139), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 key_mem_reg_6__63_ (.Q(key_mem[575]), 
	.D(FE_PHN2569_n1700), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_9__63_ (.Q(key_mem[191]), 
	.D(FE_PHN2482_n2072), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 key_mem_reg_6__31_ (.Q(key_mem[543]), 
	.D(FE_PHN2044_n1732), 
	.CK(clk_48Mhz__L6_N47));
   DFFHQX1 key_mem_reg_9__31_ (.Q(key_mem[159]), 
	.D(FE_PHN2047_n2104), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_7__110_ (.Q(key_mem[494]), 
	.D(FE_PHN2398_n1781), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_7__109_ (.Q(key_mem[493]), 
	.D(FE_PHN1045_n1782), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_7__106_ (.Q(key_mem[490]), 
	.D(FE_PHN2232_n1785), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_7__104_ (.Q(key_mem[488]), 
	.D(FE_PHN2236_n1787), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_7__112_ (.Q(key_mem[496]), 
	.D(FE_PHN1041_n1808), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_7__111_ (.Q(key_mem[495]), 
	.D(FE_PHN2536_n1809), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_7__10_ (.Q(key_mem[394]), 
	.D(FE_PHN2332_n1811), 
	.CK(clk_48Mhz__L6_N21));
   DFFHQX1 key_mem_reg_7__8_ (.Q(key_mem[392]), 
	.D(FE_PHN2622_n1813), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_7__0_ (.Q(key_mem[384]), 
	.D(FE_PHN2429_n1821), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_7__96_ (.Q(key_mem[480]), 
	.D(FE_PHN2538_n1824), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_7__80_ (.Q(key_mem[464]), 
	.D(FE_PHN2207_n1840), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_7__79_ (.Q(key_mem[463]), 
	.D(FE_PHN2494_n1841), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_7__78_ (.Q(key_mem[462]), 
	.D(FE_PHN2486_n1842), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_7__77_ (.Q(key_mem[461]), 
	.D(FE_PHN4335_n1843), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_7__74_ (.Q(key_mem[458]), 
	.D(FE_PHN2134_n1846), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_7__72_ (.Q(key_mem[456]), 
	.D(FE_PHN2148_n1848), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_7__64_ (.Q(key_mem[448]), 
	.D(FE_PHN2746_n1856), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_7__48_ (.Q(key_mem[432]), 
	.D(FE_PHN2679_n1872), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_7__47_ (.Q(key_mem[431]), 
	.D(FE_PHN2078_n1873), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_7__46_ (.Q(key_mem[430]), 
	.D(FE_PHN2543_n1874), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_7__45_ (.Q(key_mem[429]), 
	.D(FE_PHN2491_n1875), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_7__42_ (.Q(key_mem[426]), 
	.D(FE_PHN2118_n1878), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_7__40_ (.Q(key_mem[424]), 
	.D(FE_PHN2110_n1880), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_7__32_ (.Q(key_mem[416]), 
	.D(FE_PHN2620_n1888), 
	.CK(clk));
   DFFHQX1 key_mem_reg_7__16_ (.Q(key_mem[400]), 
	.D(FE_PHN2158_n1904), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_7__15_ (.Q(key_mem[399]), 
	.D(FE_PHN2189_n1905), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_7__14_ (.Q(key_mem[398]), 
	.D(FE_PHN2303_n1906), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_7__13_ (.Q(key_mem[397]), 
	.D(FE_PHN2277_n1907), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_4__112_ (.Q(key_mem[880]), 
	.D(FE_PHN2091_n1407), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_4__111_ (.Q(key_mem[879]), 
	.D(FE_PHN2654_n1408), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_4__110_ (.Q(key_mem[878]), 
	.D(FE_PHN2298_n1409), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_4__109_ (.Q(key_mem[877]), 
	.D(FE_PHN2389_n1410), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_4__106_ (.Q(key_mem[874]), 
	.D(FE_PHN1508_n1413), 
	.CK(clk_48Mhz__L6_N21));
   DFFHQX1 key_mem_reg_4__104_ (.Q(key_mem[872]), 
	.D(FE_PHN2297_n1415), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_4__16_ (.Q(key_mem[784]), 
	.D(FE_PHN2444_n1433), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_4__15_ (.Q(key_mem[783]), 
	.D(FE_PHN2441_n1434), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_4__14_ (.Q(key_mem[782]), 
	.D(FE_PHN2578_n1435), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_4__13_ (.Q(key_mem[781]), 
	.D(FE_PHN2302_n1436), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_4__10_ (.Q(key_mem[778]), 
	.D(FE_PHN626_n1439), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_4__8_ (.Q(key_mem[776]), 
	.D(FE_PHN2296_n1441), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_4__0_ (.Q(key_mem[768]), 
	.D(FE_PHN2571_n1449), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 key_mem_reg_4__96_ (.Q(key_mem[864]), 
	.D(FE_PHN2124_n1452), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_4__80_ (.Q(key_mem[848]), 
	.D(FE_PHN2717_n1468), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_4__79_ (.Q(key_mem[847]), 
	.D(FE_PHN2300_n1469), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_4__78_ (.Q(key_mem[846]), 
	.D(n1470), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_4__77_ (.Q(key_mem[845]), 
	.D(FE_PHN2558_n1471), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_4__74_ (.Q(key_mem[842]), 
	.D(FE_PHN2384_n1474), 
	.CK(clk));
   DFFHQX1 key_mem_reg_4__72_ (.Q(key_mem[840]), 
	.D(FE_PHN3965_n1476), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_4__64_ (.Q(key_mem[832]), 
	.D(FE_PHN2399_n1484), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_4__48_ (.Q(key_mem[816]), 
	.D(FE_PHN2544_n1500), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_4__47_ (.Q(key_mem[815]), 
	.D(FE_PHN4836_n1501), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_4__46_ (.Q(key_mem[814]), 
	.D(FE_PHN2376_n1502), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_4__45_ (.Q(key_mem[813]), 
	.D(FE_PHN2264_n1503), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_4__42_ (.Q(key_mem[810]), 
	.D(FE_PHN2273_n1506), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_4__40_ (.Q(key_mem[808]), 
	.D(FE_PHN2274_n1508), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_4__32_ (.Q(key_mem[800]), 
	.D(FE_PHN2648_n1516), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_10__112_ (.Q(key_mem[112]), 
	.D(FE_PHN2697_n2180), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_10__111_ (.Q(key_mem[111]), 
	.D(FE_PHN2161_n2181), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_10__110_ (.Q(key_mem[110]), 
	.D(FE_PHN2608_n2182), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_10__109_ (.Q(key_mem[109]), 
	.D(FE_PHN1527_n2183), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_10__106_ (.Q(key_mem[106]), 
	.D(FE_PHN2275_n2186), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_10__104_ (.Q(key_mem[104]), 
	.D(FE_PHN2756_n2188), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_10__96_ (.Q(key_mem[96]), 
	.D(FE_PHN2126_n2196), 
	.CK(clk));
   DFFHQX1 key_mem_reg_10__80_ (.Q(key_mem[80]), 
	.D(FE_PHN2178_n2212), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_10__79_ (.Q(key_mem[79]), 
	.D(FE_PHN2328_n2213), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_10__78_ (.Q(key_mem[78]), 
	.D(FE_PHN2083_n2214), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_10__77_ (.Q(key_mem[77]), 
	.D(FE_PHN2093_n2215), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_10__74_ (.Q(key_mem[74]), 
	.D(FE_PHN2123_n2218), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_10__72_ (.Q(key_mem[72]), 
	.D(FE_PHN2241_n2220), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_10__64_ (.Q(key_mem[64]), 
	.D(FE_PHN4452_n2228), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_10__48_ (.Q(key_mem[48]), 
	.D(FE_PHN2316_n2244), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_10__47_ (.Q(key_mem[47]), 
	.D(FE_PHN2363_n2245), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_10__46_ (.Q(key_mem[46]), 
	.D(FE_PHN2064_n2246), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_10__45_ (.Q(key_mem[45]), 
	.D(FE_PHN2257_n2247), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_10__42_ (.Q(key_mem[42]), 
	.D(FE_PHN2216_n2250), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_10__40_ (.Q(key_mem[40]), 
	.D(FE_PHN2351_n2252), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_10__32_ (.Q(key_mem[32]), 
	.D(FE_PHN2215_n2260), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_10__16_ (.Q(key_mem[16]), 
	.D(FE_PHN2415_n2276), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_10__15_ (.Q(key_mem[15]), 
	.D(FE_PHN2499_n2277), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_10__14_ (.Q(key_mem[14]), 
	.D(FE_PHN2357_n2278), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_10__13_ (.Q(key_mem[13]), 
	.D(FE_PHN1227_n2279), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_10__10_ (.Q(key_mem[10]), 
	.D(FE_PHN2182_n2282), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_10__8_ (.Q(key_mem[8]), 
	.D(FE_PHN2088_n2284), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_10__0_ (.Q(key_mem[0]), 
	.D(FE_PHN2304_n2292), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 key_mem_reg_4__122_ (.Q(key_mem[890]), 
	.D(FE_PHN2141_n1397), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_7__122_ (.Q(key_mem[506]), 
	.D(FE_PHN2373_n1798), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_10__122_ (.Q(key_mem[122]), 
	.D(FE_PHN1608_n2170), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_4__90_ (.Q(key_mem[858]), 
	.D(FE_PHN2380_n1458), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_7__90_ (.Q(key_mem[474]), 
	.D(FE_PHN2419_n1830), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_10__90_ (.Q(key_mem[90]), 
	.D(FE_PHN2279_n2202), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_4__58_ (.Q(key_mem[826]), 
	.D(FE_PHN2060_n1490), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_7__58_ (.Q(key_mem[442]), 
	.D(FE_PHN2250_n1862), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_10__58_ (.Q(key_mem[58]), 
	.D(FE_PHN2636_n2234), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_4__26_ (.Q(key_mem[794]), 
	.D(FE_PHN2625_n1522), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_7__26_ (.Q(key_mem[410]), 
	.D(FE_PHN2125_n1894), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_10__26_ (.Q(key_mem[26]), 
	.D(FE_PHN1468_n2266), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_4__125_ (.Q(key_mem[893]), 
	.D(FE_PHN2077_n1423), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_7__125_ (.Q(key_mem[509]), 
	.D(FE_PHN2467_n1795), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_10__125_ (.Q(key_mem[125]), 
	.D(FE_PHN2381_n2167), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_4__93_ (.Q(key_mem[861]), 
	.D(FE_PHN2592_n1455), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 key_mem_reg_7__93_ (.Q(key_mem[477]), 
	.D(FE_PHN2173_n1827), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_10__93_ (.Q(key_mem[93]), 
	.D(FE_PHN2058_n2199), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_4__61_ (.Q(key_mem[829]), 
	.D(FE_PHN2103_n1487), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 key_mem_reg_7__61_ (.Q(key_mem[445]), 
	.D(FE_PHN2607_n1859), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_10__61_ (.Q(key_mem[61]), 
	.D(FE_PHN2209_n2231), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_4__29_ (.Q(key_mem[797]), 
	.D(FE_PHN2416_n1519), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_7__29_ (.Q(key_mem[413]), 
	.D(FE_PHN2097_n1891), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_10__29_ (.Q(key_mem[29]), 
	.D(FE_PHN1489_n2263), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_4__126_ (.Q(key_mem[894]), 
	.D(FE_PHN2098_n1422), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_7__126_ (.Q(key_mem[510]), 
	.D(FE_PHN2336_n1794), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_10__126_ (.Q(key_mem[126]), 
	.D(FE_PHN2566_n2166), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_4__94_ (.Q(key_mem[862]), 
	.D(FE_PHN2290_n1454), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_7__94_ (.Q(key_mem[478]), 
	.D(FE_PHN2117_n1826), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_10__94_ (.Q(key_mem[94]), 
	.D(FE_PHN2086_n2198), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_4__62_ (.Q(key_mem[830]), 
	.D(FE_PHN2121_n1486), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_7__62_ (.Q(key_mem[446]), 
	.D(FE_PHN2428_n1858), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_10__62_ (.Q(key_mem[62]), 
	.D(FE_PHN2500_n2230), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_4__30_ (.Q(key_mem[798]), 
	.D(FE_PHN2591_n1518), 
	.CK(clk_48Mhz__L6_N47));
   DFFHQX1 key_mem_reg_7__30_ (.Q(key_mem[414]), 
	.D(FE_PHN2271_n1890), 
	.CK(clk_48Mhz__L6_N47));
   DFFHQX1 key_mem_reg_10__30_ (.Q(key_mem[30]), 
	.D(FE_PHN2466_n2262), 
	.CK(clk_48Mhz__L6_N47));
   DFFHQX1 key_mem_reg_4__120_ (.Q(key_mem[888]), 
	.D(FE_PHN2288_n1399), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_7__120_ (.Q(key_mem[504]), 
	.D(FE_PHN1539_n1800), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_10__120_ (.Q(key_mem[120]), 
	.D(FE_PHN1674_n2172), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_4__88_ (.Q(key_mem[856]), 
	.D(FE_PHN2531_n1460), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 key_mem_reg_7__88_ (.Q(key_mem[472]), 
	.D(FE_PHN2210_n1832), 
	.CK(clk_48Mhz__L6_N23));
   DFFHQX1 key_mem_reg_10__88_ (.Q(key_mem[88]), 
	.D(FE_PHN2147_n2204), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 key_mem_reg_4__56_ (.Q(key_mem[824]), 
	.D(FE_PHN2205_n1492), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_7__56_ (.Q(key_mem[440]), 
	.D(FE_PHN2171_n1864), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_10__56_ (.Q(key_mem[56]), 
	.D(FE_PHN2412_n2236), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_4__24_ (.Q(key_mem[792]), 
	.D(FE_PHN2478_n1524), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_7__24_ (.Q(key_mem[408]), 
	.D(FE_PHN1685_n1896), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_10__24_ (.Q(key_mem[24]), 
	.D(FE_PHN2319_n2268), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_4__127_ (.Q(key_mem[895]), 
	.D(FE_PHN2364_n1421), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_7__127_ (.Q(key_mem[511]), 
	.D(FE_PHN2596_n1793), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_10__127_ (.Q(key_mem[127]), 
	.D(FE_PHN2231_n2165), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_4__95_ (.Q(key_mem[863]), 
	.D(FE_PHN2327_n1453), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 key_mem_reg_7__95_ (.Q(key_mem[479]), 
	.D(FE_PHN2136_n1825), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_10__95_ (.Q(key_mem[95]), 
	.D(FE_PHN2186_n2197), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 key_mem_reg_4__63_ (.Q(key_mem[831]), 
	.D(FE_PHN2532_n1485), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 key_mem_reg_7__63_ (.Q(key_mem[447]), 
	.D(FE_PHN2462_n1857), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_10__63_ (.Q(key_mem[63]), 
	.D(FE_PHN2753_n2229), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 key_mem_reg_4__31_ (.Q(key_mem[799]), 
	.D(FE_PHN2618_n1517), 
	.CK(clk_48Mhz__L6_N47));
   DFFHQX1 key_mem_reg_7__31_ (.Q(key_mem[415]), 
	.D(FE_PHN2234_n1889), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_10__31_ (.Q(key_mem[31]), 
	.D(FE_PHN2193_n2261), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_8__112_ (.Q(key_mem[368]), 
	.D(FE_PHN4621_n1924), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_8__111_ (.Q(key_mem[367]), 
	.D(FE_PHN4490_n1925), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_8__110_ (.Q(key_mem[366]), 
	.D(FE_PHN4289_n1926), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_8__109_ (.Q(key_mem[365]), 
	.D(FE_PHN4444_n1927), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_8__106_ (.Q(key_mem[362]), 
	.D(FE_PHN4270_n1930), 
	.CK(clk_48Mhz__L6_N14));
   DFFHQX1 key_mem_reg_8__104_ (.Q(key_mem[360]), 
	.D(FE_PHN4941_n1932), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_8__40_ (.Q(key_mem[296]), 
	.D(FE_PHN4338_n1938), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_8__32_ (.Q(key_mem[288]), 
	.D(FE_PHN4339_n1946), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_8__16_ (.Q(key_mem[272]), 
	.D(FE_PHN4821_n1962), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_8__15_ (.Q(key_mem[271]), 
	.D(FE_PHN4278_n1963), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_8__14_ (.Q(key_mem[270]), 
	.D(FE_PHN4345_n1964), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_8__13_ (.Q(key_mem[269]), 
	.D(FE_PHN4877_n1965), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_8__10_ (.Q(key_mem[266]), 
	.D(FE_PHN4312_n1968), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_8__8_ (.Q(key_mem[264]), 
	.D(FE_PHN4585_n1970), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_8__0_ (.Q(key_mem[256]), 
	.D(FE_PHN4953_n1978), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_8__96_ (.Q(key_mem[352]), 
	.D(FE_PHN4985_n1981), 
	.CK(clk));
   DFFHQX1 key_mem_reg_8__80_ (.Q(key_mem[336]), 
	.D(FE_PHN4065_n1997), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_8__79_ (.Q(key_mem[335]), 
	.D(FE_PHN3856_n1998), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_8__78_ (.Q(key_mem[334]), 
	.D(FE_PHN4918_n1999), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_8__77_ (.Q(key_mem[333]), 
	.D(FE_PHN4053_n2000), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_8__74_ (.Q(key_mem[330]), 
	.D(FE_PHN4075_n2003), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_8__72_ (.Q(key_mem[328]), 
	.D(FE_PHN4572_n2005), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_8__64_ (.Q(key_mem[320]), 
	.D(FE_PHN4305_n2013), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_8__48_ (.Q(key_mem[304]), 
	.D(FE_PHN4299_n2029), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_8__47_ (.Q(key_mem[303]), 
	.D(FE_PHN4689_n2030), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_8__46_ (.Q(key_mem[302]), 
	.D(FE_PHN4712_n2031), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_8__45_ (.Q(key_mem[301]), 
	.D(FE_PHN4258_n2032), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_8__42_ (.Q(key_mem[298]), 
	.D(FE_PHN4849_n2035), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_5__112_ (.Q(key_mem[752]), 
	.D(FE_PHN4426_n1540), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_5__111_ (.Q(key_mem[751]), 
	.D(FE_PHN4183_n1541), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_5__110_ (.Q(key_mem[750]), 
	.D(FE_PHN4061_n1542), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_5__109_ (.Q(key_mem[749]), 
	.D(FE_PHN4592_n1543), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_5__106_ (.Q(key_mem[746]), 
	.D(FE_PHN1576_n1546), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_5__104_ (.Q(key_mem[744]), 
	.D(FE_PHN4602_n1548), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_5__48_ (.Q(key_mem[688]), 
	.D(FE_PHN4964_n1558), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_5__47_ (.Q(key_mem[687]), 
	.D(FE_PHN4550_n1559), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_5__46_ (.Q(key_mem[686]), 
	.D(FE_PHN4349_n1560), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_5__45_ (.Q(key_mem[685]), 
	.D(FE_PHN4797_n1561), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_5__42_ (.Q(key_mem[682]), 
	.D(FE_PHN4760_n1564), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_5__40_ (.Q(key_mem[680]), 
	.D(FE_PHN4651_n1566), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_5__32_ (.Q(key_mem[672]), 
	.D(FE_PHN4231_n1574), 
	.CK(clk));
   DFFHQX1 key_mem_reg_5__16_ (.Q(key_mem[656]), 
	.D(FE_PHN4219_n1590), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_5__15_ (.Q(key_mem[655]), 
	.D(FE_PHN4291_n1591), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_5__14_ (.Q(key_mem[654]), 
	.D(FE_PHN4469_n1592), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_5__13_ (.Q(key_mem[653]), 
	.D(FE_PHN1585_n1593), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_5__10_ (.Q(key_mem[650]), 
	.D(FE_PHN1736_n1596), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_5__8_ (.Q(key_mem[648]), 
	.D(FE_PHN4864_n1598), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_5__0_ (.Q(key_mem[640]), 
	.D(FE_PHN4093_n1606), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_5__96_ (.Q(key_mem[736]), 
	.D(FE_PHN4225_n1609), 
	.CK(clk));
   DFFHQX1 key_mem_reg_5__80_ (.Q(key_mem[720]), 
	.D(FE_PHN4436_n1625), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_5__79_ (.Q(key_mem[719]), 
	.D(FE_PHN4082_n1626), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_5__78_ (.Q(key_mem[718]), 
	.D(FE_PHN4098_n1627), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_5__77_ (.Q(key_mem[717]), 
	.D(FE_PHN4463_n1628), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_5__74_ (.Q(key_mem[714]), 
	.D(FE_PHN3855_n1631), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_5__72_ (.Q(key_mem[712]), 
	.D(FE_PHN4326_n1633), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_5__64_ (.Q(key_mem[704]), 
	.D(FE_PHN4690_n1641), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_5__121_ (.Q(key_mem[761]), 
	.D(FE_PHN1654_n1531), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_8__121_ (.Q(key_mem[377]), 
	.D(FE_PHN4632_n1915), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_5__89_ (.Q(key_mem[729]), 
	.D(FE_PHN4100_n1616), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_8__89_ (.Q(key_mem[345]), 
	.D(FE_PHN4480_n1988), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_5__57_ (.Q(key_mem[697]), 
	.D(FE_PHN4313_n1648), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_8__57_ (.Q(key_mem[313]), 
	.D(FE_PHN4348_n2020), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_5__25_ (.Q(key_mem[665]), 
	.D(FE_PHN1676_n1581), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_8__25_ (.Q(key_mem[281]), 
	.D(FE_PHN4365_n1953), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_5__122_ (.Q(key_mem[762]), 
	.D(FE_PHN4387_n1530), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_8__122_ (.Q(key_mem[378]), 
	.D(FE_PHN4571_n1914), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_5__90_ (.Q(key_mem[730]), 
	.D(FE_PHN4768_n1615), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_8__90_ (.Q(key_mem[346]), 
	.D(FE_PHN4779_n1987), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_5__58_ (.Q(key_mem[698]), 
	.D(FE_PHN4844_n1647), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_8__58_ (.Q(key_mem[314]), 
	.D(FE_PHN4609_n2019), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_5__26_ (.Q(key_mem[666]), 
	.D(FE_PHN1611_n1580), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_8__26_ (.Q(key_mem[282]), 
	.D(FE_PHN4566_n1952), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_5__123_ (.Q(key_mem[763]), 
	.D(FE_PHN4771_n1529), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_8__123_ (.Q(key_mem[379]), 
	.D(FE_PHN3951_n1913), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_5__91_ (.Q(key_mem[731]), 
	.D(FE_PHN4830_n1614), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_8__91_ (.Q(key_mem[347]), 
	.D(FE_PHN4584_n1986), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_5__59_ (.Q(key_mem[699]), 
	.D(FE_PHN4044_n1646), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_8__59_ (.Q(key_mem[315]), 
	.D(FE_PHN4375_n2018), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_5__27_ (.Q(key_mem[667]), 
	.D(FE_PHN1796_n1579), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_8__27_ (.Q(key_mem[283]), 
	.D(FE_PHN4092_n1951), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_5__124_ (.Q(key_mem[764]), 
	.D(FE_PHN4685_n1528), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_8__124_ (.Q(key_mem[380]), 
	.D(FE_PHN4788_n1912), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_5__92_ (.Q(key_mem[732]), 
	.D(FE_PHN4635_n1613), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_8__92_ (.Q(key_mem[348]), 
	.D(FE_PHN4518_n1985), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_5__60_ (.Q(key_mem[700]), 
	.D(FE_PHN4474_n1645), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 key_mem_reg_8__60_ (.Q(key_mem[316]), 
	.D(FE_PHN4883_n2017), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_5__28_ (.Q(key_mem[668]), 
	.D(FE_PHN1693_n1578), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_8__28_ (.Q(key_mem[284]), 
	.D(FE_PHN4497_n1950), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_5__125_ (.Q(key_mem[765]), 
	.D(FE_PHN4704_n1527), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_8__125_ (.Q(key_mem[381]), 
	.D(FE_PHN4255_n1911), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_5__93_ (.Q(key_mem[733]), 
	.D(FE_PHN4950_n1612), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_8__93_ (.Q(key_mem[349]), 
	.D(FE_PHN4894_n1984), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 key_mem_reg_5__61_ (.Q(key_mem[701]), 
	.D(FE_PHN4377_n1644), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_8__61_ (.Q(key_mem[317]), 
	.D(FE_PHN4659_n2016), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_5__29_ (.Q(key_mem[669]), 
	.D(FE_PHN1570_n1577), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_8__29_ (.Q(key_mem[285]), 
	.D(FE_PHN4695_n1949), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_5__126_ (.Q(key_mem[766]), 
	.D(FE_PHN4863_n1526), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_8__126_ (.Q(key_mem[382]), 
	.D(FE_PHN4488_n1910), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_5__94_ (.Q(key_mem[734]), 
	.D(FE_PHN4802_n1611), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_8__94_ (.Q(key_mem[350]), 
	.D(FE_PHN4264_n1983), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_5__62_ (.Q(key_mem[702]), 
	.D(FE_PHN4792_n1643), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_8__62_ (.Q(key_mem[318]), 
	.D(FE_PHN4795_n2015), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_5__30_ (.Q(key_mem[670]), 
	.D(FE_PHN3949_n1576), 
	.CK(clk_48Mhz__L6_N47));
   DFFHQX1 key_mem_reg_8__30_ (.Q(key_mem[286]), 
	.D(FE_PHN3979_n1948), 
	.CK(clk_48Mhz__L6_N47));
   DFFHQX1 key_mem_reg_5__120_ (.Q(key_mem[760]), 
	.D(FE_PHN4644_n1532), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_8__120_ (.Q(key_mem[376]), 
	.D(FE_PHN4987_n1916), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_5__88_ (.Q(key_mem[728]), 
	.D(FE_PHN4832_n1617), 
	.CK(clk_48Mhz__L6_N23));
   DFFHQX1 key_mem_reg_8__88_ (.Q(key_mem[344]), 
	.D(FE_PHN4875_n1989), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 key_mem_reg_5__56_ (.Q(key_mem[696]), 
	.D(FE_PHN4852_n1649), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_8__56_ (.Q(key_mem[312]), 
	.D(FE_PHN4088_n2021), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_5__24_ (.Q(key_mem[664]), 
	.D(FE_PHN4598_n1582), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_8__24_ (.Q(key_mem[280]), 
	.D(FE_PHN4245_n1954), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_5__127_ (.Q(key_mem[767]), 
	.D(FE_PHN4611_n1525), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_8__127_ (.Q(key_mem[383]), 
	.D(FE_PHN4243_n1909), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_5__95_ (.Q(key_mem[735]), 
	.D(FE_PHN4654_n1610), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_8__95_ (.Q(key_mem[351]), 
	.D(FE_PHN4582_n1982), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 key_mem_reg_5__63_ (.Q(key_mem[703]), 
	.D(FE_PHN4737_n1642), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_8__63_ (.Q(key_mem[319]), 
	.D(FE_PHN4617_n2014), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 key_mem_reg_5__31_ (.Q(key_mem[671]), 
	.D(FE_PHN4630_n1575), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_8__31_ (.Q(key_mem[287]), 
	.D(FE_PHN4558_n1947), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 prev_key1_reg_reg_55_ (.Q(prev_key1_reg[55]), 
	.D(FE_PHN4899_n2365), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 prev_key1_reg_reg_54_ (.Q(prev_key1_reg[54]), 
	.D(FE_PHN4809_n2366), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 prev_key1_reg_reg_53_ (.Q(prev_key1_reg[53]), 
	.D(FE_PHN4189_n2367), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 prev_key1_reg_reg_52_ (.Q(prev_key1_reg[52]), 
	.D(FE_PHN4629_n2368), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 prev_key1_reg_reg_51_ (.Q(prev_key1_reg[51]), 
	.D(FE_PHN4767_n2369), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 prev_key1_reg_reg_50_ (.Q(prev_key1_reg[50]), 
	.D(FE_PHN4940_n2370), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 prev_key1_reg_reg_49_ (.Q(prev_key1_reg[49]), 
	.D(FE_PHN4851_n2371), 
	.CK(clk_48Mhz__L6_N11));
   DFFHQX1 prev_key1_reg_reg_48_ (.Q(prev_key1_reg[48]), 
	.D(FE_PHN715_n2372), 
	.CK(clk_48Mhz__L6_N11));
   DFFHQX1 prev_key1_reg_reg_47_ (.Q(prev_key1_reg[47]), 
	.D(FE_PHN1315_n2373), 
	.CK(clk_48Mhz__L6_N9));
   DFFHQX1 prev_key1_reg_reg_46_ (.Q(prev_key1_reg[46]), 
	.D(FE_PHN714_n2374), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 prev_key1_reg_reg_45_ (.Q(prev_key1_reg[45]), 
	.D(FE_PHN4703_n2375), 
	.CK(clk_48Mhz__L6_N27));
   DFFHQX1 prev_key1_reg_reg_44_ (.Q(prev_key1_reg[44]), 
	.D(FE_PHN4954_n2376), 
	.CK(clk_48Mhz__L6_N27));
   DFFHQX1 prev_key1_reg_reg_43_ (.Q(prev_key1_reg[43]), 
	.D(FE_PHN4118_n2377), 
	.CK(clk_48Mhz__L6_N23));
   DFFHQX1 prev_key1_reg_reg_42_ (.Q(prev_key1_reg[42]), 
	.D(FE_PHN4417_n2378), 
	.CK(clk_48Mhz__L6_N14));
   DFFHQX1 prev_key1_reg_reg_41_ (.Q(prev_key1_reg[41]), 
	.D(FE_PHN4948_n2379), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 prev_key1_reg_reg_40_ (.Q(prev_key1_reg[40]), 
	.D(FE_PHN4285_n2380), 
	.CK(clk_48Mhz__L6_N11));
   DFFHQX1 prev_key1_reg_reg_39_ (.Q(prev_key1_reg[39]), 
	.D(FE_PHN1312_n2381), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 prev_key1_reg_reg_38_ (.Q(prev_key1_reg[38]), 
	.D(FE_PHN4462_n2382), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 prev_key1_reg_reg_37_ (.Q(prev_key1_reg[37]), 
	.D(FE_PHN4783_n2383), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 prev_key1_reg_reg_36_ (.Q(prev_key1_reg[36]), 
	.D(FE_PHN4564_n2384), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 prev_key1_reg_reg_35_ (.Q(prev_key1_reg[35]), 
	.D(FE_PHN4942_n2385), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 prev_key1_reg_reg_34_ (.Q(prev_key1_reg[34]), 
	.D(FE_PHN4027_n2386), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 prev_key1_reg_reg_33_ (.Q(prev_key1_reg[33]), 
	.D(FE_PHN4396_n2387), 
	.CK(clk));
   DFFHQX1 prev_key1_reg_reg_32_ (.Q(prev_key1_reg[32]), 
	.D(FE_PHN4530_n2388), 
	.CK(clk));
   DFFHQX1 prev_key1_reg_reg_119_ (.Q(prev_key1_reg[119]), 
	.D(FE_PHN4477_n2301), 
	.CK(clk_48Mhz__L6_N9));
   DFFHQX1 prev_key1_reg_reg_118_ (.Q(prev_key1_reg[118]), 
	.D(FE_PHN4812_n2302), 
	.CK(clk_48Mhz__L6_N10));
   DFFHQX1 prev_key1_reg_reg_117_ (.Q(prev_key1_reg[117]), 
	.D(FE_PHN4117_n2303), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 prev_key1_reg_reg_116_ (.Q(prev_key1_reg[116]), 
	.D(FE_PHN4973_n2304), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 prev_key1_reg_reg_115_ (.Q(prev_key1_reg[115]), 
	.D(FE_PHN4658_n2305), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 prev_key1_reg_reg_114_ (.Q(prev_key1_reg[114]), 
	.D(FE_PHN4412_n2306), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 prev_key1_reg_reg_113_ (.Q(prev_key1_reg[113]), 
	.D(FE_PHN4536_n2307), 
	.CK(clk_48Mhz__L6_N11));
   DFFHQX1 prev_key1_reg_reg_112_ (.Q(prev_key1_reg[112]), 
	.D(FE_PHN4814_n2308), 
	.CK(clk_48Mhz__L6_N11));
   DFFHQX1 prev_key1_reg_reg_111_ (.Q(prev_key1_reg[111]), 
	.D(FE_PHN4575_n2309), 
	.CK(clk_48Mhz__L6_N9));
   DFFHQX1 prev_key1_reg_reg_110_ (.Q(prev_key1_reg[110]), 
	.D(FE_PHN4591_n2310), 
	.CK(clk_48Mhz__L6_N9));
   DFFHQX1 prev_key1_reg_reg_109_ (.Q(prev_key1_reg[109]), 
	.D(FE_PHN4489_n2311), 
	.CK(clk_48Mhz__L6_N14));
   DFFHQX1 prev_key1_reg_reg_108_ (.Q(prev_key1_reg[108]), 
	.D(FE_PHN4968_n2312), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 prev_key1_reg_reg_107_ (.Q(prev_key1_reg[107]), 
	.D(FE_PHN4884_n2313), 
	.CK(clk_48Mhz__L6_N14));
   DFFHQX1 prev_key1_reg_reg_106_ (.Q(prev_key1_reg[106]), 
	.D(FE_PHN4787_n2314), 
	.CK(clk_48Mhz__L6_N14));
   DFFHQX1 prev_key1_reg_reg_105_ (.Q(prev_key1_reg[105]), 
	.D(FE_PHN4845_n2315), 
	.CK(clk_48Mhz__L6_N11));
   DFFHQX1 prev_key1_reg_reg_104_ (.Q(prev_key1_reg[104]), 
	.D(FE_PHN4650_n2316), 
	.CK(clk_48Mhz__L6_N6));
   DFFHQX1 prev_key1_reg_reg_103_ (.Q(prev_key1_reg[103]), 
	.D(FE_PHN4333_n2317), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 prev_key1_reg_reg_102_ (.Q(prev_key1_reg[102]), 
	.D(FE_PHN4195_n2318), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 prev_key1_reg_reg_101_ (.Q(prev_key1_reg[101]), 
	.D(FE_PHN4876_n2319), 
	.CK(clk_48Mhz__L6_N23));
   DFFHQX1 prev_key1_reg_reg_100_ (.Q(prev_key1_reg[100]), 
	.D(FE_PHN4715_n2320), 
	.CK(clk_48Mhz__L6_N23));
   DFFHQX1 prev_key1_reg_reg_99_ (.Q(prev_key1_reg[99]), 
	.D(FE_PHN4397_n2321), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 prev_key1_reg_reg_98_ (.Q(prev_key1_reg[98]), 
	.D(FE_PHN4457_n2322), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 prev_key1_reg_reg_97_ (.Q(prev_key1_reg[97]), 
	.D(FE_PHN4269_n2323), 
	.CK(clk));
   DFFHQX1 prev_key1_reg_reg_96_ (.Q(prev_key1_reg[96]), 
	.D(FE_PHN4664_n2324), 
	.CK(clk));
   DFFHQX1 prev_key1_reg_reg_89_ (.Q(prev_key1_reg[89]), 
	.D(FE_PHN4097_n2331), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 prev_key1_reg_reg_90_ (.Q(prev_key1_reg[90]), 
	.D(FE_PHN4673_n2330), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 prev_key1_reg_reg_91_ (.Q(prev_key1_reg[91]), 
	.D(FE_PHN4263_n2329), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 prev_key1_reg_reg_92_ (.Q(prev_key1_reg[92]), 
	.D(FE_PHN4304_n2328), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 prev_key1_reg_reg_93_ (.Q(prev_key1_reg[93]), 
	.D(FE_PHN4888_n2327), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 prev_key1_reg_reg_94_ (.Q(prev_key1_reg[94]), 
	.D(FE_PHN4874_n2326), 
	.CK(clk_48Mhz__L6_N6));
   DFFHQX1 prev_key1_reg_reg_88_ (.Q(prev_key1_reg[88]), 
	.D(FE_PHN4840_n2332), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 prev_key1_reg_reg_95_ (.Q(prev_key1_reg[95]), 
	.D(FE_PHN4448_n2325), 
	.CK(clk_48Mhz__L6_N9));
   DFFHQX1 prev_key1_reg_reg_57_ (.Q(prev_key1_reg[57]), 
	.D(FE_PHN5028_n2363), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 prev_key1_reg_reg_58_ (.Q(prev_key1_reg[58]), 
	.D(FE_PHN5017_n2362), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 prev_key1_reg_reg_59_ (.Q(prev_key1_reg[59]), 
	.D(FE_PHN5009_n2361), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 prev_key1_reg_reg_60_ (.Q(prev_key1_reg[60]), 
	.D(FE_PHN5015_n2360), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 prev_key1_reg_reg_61_ (.Q(prev_key1_reg[61]), 
	.D(FE_PHN5036_n2359), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 prev_key1_reg_reg_62_ (.Q(prev_key1_reg[62]), 
	.D(FE_PHN4994_n2358), 
	.CK(clk_48Mhz__L6_N6));
   DFFHQX1 prev_key1_reg_reg_56_ (.Q(prev_key1_reg[56]), 
	.D(FE_PHN747_n2364), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 prev_key1_reg_reg_63_ (.Q(prev_key1_reg[63]), 
	.D(FE_PHN5010_n2357), 
	.CK(clk_48Mhz__L6_N6));
   DFFHQX1 prev_key1_reg_reg_121_ (.Q(prev_key1_reg[121]), 
	.D(FE_PHN4992_n2299), 
	.CK(clk_48Mhz__L6_N8));
   DFFHQX1 prev_key1_reg_reg_122_ (.Q(prev_key1_reg[122]), 
	.D(FE_PHN4986_n2298), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 prev_key1_reg_reg_123_ (.Q(prev_key1_reg[123]), 
	.D(FE_PHN5021_n2297), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 prev_key1_reg_reg_124_ (.Q(prev_key1_reg[124]), 
	.D(FE_PHN5005_n2296), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 prev_key1_reg_reg_125_ (.Q(prev_key1_reg[125]), 
	.D(FE_PHN5014_n2295), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 prev_key1_reg_reg_126_ (.Q(prev_key1_reg[126]), 
	.D(FE_PHN1211_n2294), 
	.CK(clk_48Mhz__L6_N6));
   DFFHQX1 prev_key1_reg_reg_120_ (.Q(prev_key1_reg[120]), 
	.D(FE_PHN5018_n2300), 
	.CK(clk_48Mhz__L6_N8));
   DFFHQX1 prev_key1_reg_reg_127_ (.Q(prev_key1_reg[127]), 
	.D(FE_PHN5023_n2293), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 key_mem_reg_3__112_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1008]), 
	.D(FE_PHN2748_n1284), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_3__111_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1007]), 
	.D(FE_PHN2584_n1285), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 key_mem_reg_3__110_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1006]), 
	.D(FE_PHN2734_n1286), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_3__109_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1005]), 
	.D(FE_PHN2567_n1287), 
	.CK(clk_48Mhz__L6_N19));
   DFFRHQX1 key_mem_reg_3__106_ (.RN(FE_OFN39_reset_n), 
	.Q(key_mem[1002]), 
	.D(FE_PHN1075_n1290), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 key_mem_reg_3__104_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1000]), 
	.D(FE_PHN2694_n1292), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 key_mem_reg_3__96_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[992]), 
	.D(FE_PHN2624_n1300), 
	.CK(clk_48Mhz__L6_N25));
   DFFRHQX1 key_mem_reg_3__80_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[976]), 
	.D(FE_PHN2594_n1316), 
	.CK(clk_48Mhz__L6_N7));
   DFFRHQX1 key_mem_reg_3__79_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[975]), 
	.D(FE_PHN806_n1317), 
	.CK(clk_48Mhz__L6_N3));
   DFFRHQX1 key_mem_reg_3__78_ (.RN(FE_OFN42_reset_n), 
	.Q(key_mem[974]), 
	.D(FE_PHN2527_n1318), 
	.CK(clk_48Mhz__L6_N1));
   DFFRHQX1 key_mem_reg_3__77_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[973]), 
	.D(FE_PHN2773_n1319), 
	.CK(clk_48Mhz__L6_N7));
   DFFRHQX1 key_mem_reg_3__74_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[970]), 
	.D(FE_PHN2656_n1322), 
	.CK(clk_48Mhz__L6_N25));
   DFFRHQX1 key_mem_reg_3__72_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[968]), 
	.D(FE_PHN2653_n1324), 
	.CK(clk_48Mhz__L6_N3));
   DFFRHQX1 key_mem_reg_3__64_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[960]), 
	.D(FE_PHN2765_n1332), 
	.CK(clk_48Mhz__L6_N25));
   DFFRHQX1 key_mem_reg_3__48_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[944]), 
	.D(FE_PHN2783_n1348), 
	.CK(clk_48Mhz__L6_N24));
   DFFRHQX1 key_mem_reg_3__47_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[943]), 
	.D(FE_PHN2726_n1349), 
	.CK(clk_48Mhz__L6_N31));
   DFFRHQX1 key_mem_reg_3__46_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[942]), 
	.D(FE_PHN2741_n1350), 
	.CK(clk_48Mhz__L6_N24));
   DFFRHQX1 key_mem_reg_3__45_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[941]), 
	.D(FE_PHN2735_n1351), 
	.CK(clk_48Mhz__L6_N33));
   DFFRHQX1 key_mem_reg_3__42_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[938]), 
	.D(FE_PHN737_n1354), 
	.CK(clk_48Mhz__L6_N31));
   DFFRHQX1 key_mem_reg_3__40_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[936]), 
	.D(FE_PHN2762_n1356), 
	.CK(clk_48Mhz__L6_N24));
   DFFRHQX1 key_mem_reg_3__32_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[928]), 
	.D(FE_PHN710_n1364), 
	.CK(clk_48Mhz__L6_N7));
   DFFRHQX1 key_mem_reg_3__16_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[912]), 
	.D(FE_PHN2764_n1380), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_3__15_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[911]), 
	.D(FE_PHN593_n1381), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_3__14_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[910]), 
	.D(FE_PHN2613_n1382), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_3__13_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[909]), 
	.D(FE_PHN2686_n1383), 
	.CK(clk_48Mhz__L6_N19));
   DFFRHQX1 key_mem_reg_3__10_ (.RN(FE_OFN55_reset_n), 
	.Q(key_mem[906]), 
	.D(FE_PHN997_n1386), 
	.CK(clk_48Mhz__L6_N22));
   DFFRHQX1 key_mem_reg_3__8_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[904]), 
	.D(FE_PHN2651_n1388), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 key_mem_reg_3__0_ (.RN(FE_OFN42_reset_n), 
	.Q(key_mem[896]), 
	.D(FE_PHN957_n1396), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 key_mem_reg_3__122_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1018]), 
	.D(FE_PHN2510_n1274), 
	.CK(clk_48Mhz__L6_N22));
   DFFRHQX1 key_mem_reg_3__90_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[986]), 
	.D(FE_PHN991_n1306), 
	.CK(clk_48Mhz__L6_N17));
   DFFRHQX1 key_mem_reg_3__58_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[954]), 
	.D(FE_PHN2768_n1338), 
	.CK(clk_48Mhz__L6_N17));
   DFFRHQX1 key_mem_reg_3__26_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[922]), 
	.D(FE_PHN2623_n1370), 
	.CK(clk_48Mhz__L6_N19));
   DFFRHQX1 key_mem_reg_3__125_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1021]), 
	.D(FE_PHN2646_n1271), 
	.CK(clk_48Mhz__L6_N12));
   DFFRHQX1 key_mem_reg_3__93_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[989]), 
	.D(FE_PHN2718_n1303), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 key_mem_reg_3__61_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[957]), 
	.D(FE_PHN722_n1335), 
	.CK(clk_48Mhz__L6_N33));
   DFFRHQX1 key_mem_reg_3__29_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[925]), 
	.D(FE_PHN2497_n1367), 
	.CK(clk_48Mhz__L6_N22));
   DFFRHQX1 key_mem_reg_3__126_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1022]), 
	.D(FE_PHN2663_n1270), 
	.CK(clk_48Mhz__L6_N42));
   DFFRHQX1 key_mem_reg_3__94_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[990]), 
	.D(FE_PHN2691_n1302), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 key_mem_reg_3__62_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[958]), 
	.D(FE_PHN2458_n1334), 
	.CK(clk_48Mhz__L6_N32));
   DFFRHQX1 key_mem_reg_3__30_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[926]), 
	.D(FE_PHN723_n1366), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_3__120_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1016]), 
	.D(FE_PHN2737_n1276), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_3__88_ (.RN(FE_OFN45_reset_n), 
	.Q(key_mem[984]), 
	.D(FE_PHN646_n1308), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 key_mem_reg_3__56_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[952]), 
	.D(FE_PHN2751_n1340), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_3__24_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[920]), 
	.D(FE_PHN2699_n1372), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_3__127_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1023]), 
	.D(FE_PHN2736_n1269), 
	.CK(clk_48Mhz__L6_N42));
   DFFRHQX1 key_mem_reg_3__95_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[991]), 
	.D(FE_PHN2724_n1301), 
	.CK(clk_48Mhz__L6_N1));
   DFFRHQX1 key_mem_reg_3__63_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[959]), 
	.D(FE_PHN2631_n1333), 
	.CK(clk_48Mhz__L6_N32));
   DFFRHQX1 key_mem_reg_3__31_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[927]), 
	.D(FE_PHN738_n1365), 
	.CK(clk_48Mhz__L6_N42));
   DFFRHQX1 key_mem_reg_2__112_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1136]), 
	.D(FE_PHN4815_n1156), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_2__111_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1135]), 
	.D(FE_PHN4765_n1157), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 key_mem_reg_2__110_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1134]), 
	.D(FE_PHN4853_n1158), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_2__109_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1133]), 
	.D(FE_PHN4738_n1159), 
	.CK(clk_48Mhz__L6_N19));
   DFFRHQX1 key_mem_reg_2__106_ (.RN(FE_OFN39_reset_n), 
	.Q(key_mem[1130]), 
	.D(FE_PHN1847_n1162), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 key_mem_reg_2__104_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1128]), 
	.D(FE_PHN4782_n1164), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 key_mem_reg_2__96_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1120]), 
	.D(FE_PHN4824_n1172), 
	.CK(clk));
   DFFRHQX1 key_mem_reg_2__80_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1104]), 
	.D(FE_PHN4646_n1188), 
	.CK(clk_48Mhz__L6_N7));
   DFFRHQX1 key_mem_reg_2__79_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1103]), 
	.D(FE_PHN4856_n1189), 
	.CK(clk_48Mhz__L6_N3));
   DFFRHQX1 key_mem_reg_2__78_ (.RN(FE_OFN42_reset_n), 
	.Q(key_mem[1102]), 
	.D(FE_PHN803_n1190), 
	.CK(clk_48Mhz__L6_N1));
   DFFRHQX1 key_mem_reg_2__77_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1101]), 
	.D(FE_PHN4961_n1191), 
	.CK(clk_48Mhz__L6_N7));
   DFFRHQX1 key_mem_reg_2__74_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1098]), 
	.D(FE_PHN4903_n1194), 
	.CK(clk));
   DFFRHQX1 key_mem_reg_2__72_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1096]), 
	.D(FE_PHN973_n1196), 
	.CK(clk_48Mhz__L6_N3));
   DFFRHQX1 key_mem_reg_2__64_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1088]), 
	.D(FE_PHN4823_n1204), 
	.CK(clk_48Mhz__L6_N28));
   DFFRHQX1 key_mem_reg_2__48_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1072]), 
	.D(FE_PHN4900_n1220), 
	.CK(clk_48Mhz__L6_N24));
   DFFRHQX1 key_mem_reg_2__47_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1071]), 
	.D(FE_PHN4892_n1221), 
	.CK(clk_48Mhz__L6_N31));
   DFFRHQX1 key_mem_reg_2__46_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1070]), 
	.D(FE_PHN4301_n1222), 
	.CK(clk_48Mhz__L6_N24));
   DFFRHQX1 key_mem_reg_2__45_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1069]), 
	.D(FE_PHN4829_n1223), 
	.CK(clk_48Mhz__L6_N31));
   DFFRHQX1 key_mem_reg_2__42_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1066]), 
	.D(FE_PHN4656_n1226), 
	.CK(clk_48Mhz__L6_N31));
   DFFRHQX1 key_mem_reg_2__40_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1064]), 
	.D(FE_PHN4843_n1228), 
	.CK(clk_48Mhz__L6_N24));
   DFFRHQX1 key_mem_reg_2__32_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1056]), 
	.D(FE_PHN728_n1236), 
	.CK(clk_48Mhz__L6_N7));
   DFFRHQX1 key_mem_reg_2__16_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1040]), 
	.D(FE_PHN4922_n1252), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_2__15_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1039]), 
	.D(FE_PHN4911_n1253), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 key_mem_reg_2__14_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1038]), 
	.D(FE_PHN959_n1254), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_2__13_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1037]), 
	.D(FE_PHN4746_n1255), 
	.CK(clk_48Mhz__L6_N19));
   DFFRHQX1 key_mem_reg_2__10_ (.RN(FE_OFN55_reset_n), 
	.Q(key_mem[1034]), 
	.D(FE_PHN1709_n1258), 
	.CK(clk_48Mhz__L6_N22));
   DFFRHQX1 key_mem_reg_2__8_ (.RN(FE_OFN45_reset_n), 
	.Q(key_mem[1032]), 
	.D(FE_PHN4438_n1260), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 key_mem_reg_2__0_ (.RN(FE_OFN42_reset_n), 
	.Q(key_mem[1024]), 
	.D(FE_PHN1022_n1268), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 key_mem_reg_2__121_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1145]), 
	.D(FE_PHN4699_n1147), 
	.CK(clk_48Mhz__L6_N18));
   DFFRHQX1 key_mem_reg_2__89_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1113]), 
	.D(FE_PHN4967_n1179), 
	.CK(clk_48Mhz__L6_N33));
   DFFRHQX1 key_mem_reg_2__57_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1081]), 
	.D(FE_PHN4583_n1211), 
	.CK(clk_48Mhz__L6_N20));
   DFFRHQX1 key_mem_reg_2__25_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1049]), 
	.D(FE_PHN4943_n1243), 
	.CK(clk_48Mhz__L6_N18));
   DFFRHQX1 key_mem_reg_2__122_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1146]), 
	.D(FE_PHN807_n1146), 
	.CK(clk_48Mhz__L6_N19));
   DFFRHQX1 key_mem_reg_2__90_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1114]), 
	.D(FE_PHN4981_n1178), 
	.CK(clk_48Mhz__L6_N17));
   DFFRHQX1 key_mem_reg_2__58_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1082]), 
	.D(FE_PHN4991_n1210), 
	.CK(clk_48Mhz__L6_N17));
   DFFRHQX1 key_mem_reg_2__26_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1050]), 
	.D(FE_PHN4425_n1242), 
	.CK(clk_48Mhz__L6_N19));
   DFFRHQX1 key_mem_reg_2__123_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1147]), 
	.D(FE_PHN4639_n1145), 
	.CK(clk_48Mhz__L6_N19));
   DFFRHQX1 key_mem_reg_2__91_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1115]), 
	.D(FE_PHN4764_n1177), 
	.CK(clk_48Mhz__L6_N26));
   DFFRHQX1 key_mem_reg_2__59_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1083]), 
	.D(FE_PHN4924_n1209), 
	.CK(clk_48Mhz__L6_N17));
   DFFRHQX1 key_mem_reg_2__27_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1051]), 
	.D(FE_PHN4811_n1241), 
	.CK(clk_48Mhz__L6_N18));
   DFFRHQX1 key_mem_reg_2__124_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1148]), 
	.D(FE_PHN4882_n1144), 
	.CK(clk_48Mhz__L6_N12));
   DFFRHQX1 key_mem_reg_2__92_ (.RN(FE_OFN43_reset_n), 
	.Q(key_mem[1116]), 
	.D(FE_PHN4605_n1176), 
	.CK(clk_48Mhz__L6_N20));
   DFFRHQX1 key_mem_reg_2__60_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1084]), 
	.D(FE_PHN4946_n1208), 
	.CK(clk_48Mhz__L6_N33));
   DFFRHQX1 key_mem_reg_2__28_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1052]), 
	.D(FE_PHN1801_n1240), 
	.CK(clk_48Mhz__L6_N22));
   DFFRHQX1 key_mem_reg_2__125_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1149]), 
	.D(FE_PHN961_n1143), 
	.CK(clk_48Mhz__L6_N12));
   DFFRHQX1 key_mem_reg_2__93_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1117]), 
	.D(FE_PHN632_n1175), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 key_mem_reg_2__61_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1085]), 
	.D(FE_PHN4982_n1207), 
	.CK(clk_48Mhz__L6_N33));
   DFFRHQX1 key_mem_reg_2__29_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1053]), 
	.D(FE_PHN4976_n1239), 
	.CK(clk_48Mhz__L6_N22));
   DFFRHQX1 key_mem_reg_2__126_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1150]), 
	.D(FE_PHN4906_n1142), 
	.CK(clk_48Mhz__L6_N42));
   DFFRHQX1 key_mem_reg_2__94_ (.RN(FE_OFN42_reset_n), 
	.Q(key_mem[1118]), 
	.D(FE_PHN4668_n1174), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 key_mem_reg_2__62_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1086]), 
	.D(FE_PHN812_n1206), 
	.CK(clk_48Mhz__L6_N32));
   DFFRHQX1 key_mem_reg_2__30_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1054]), 
	.D(FE_PHN4337_n1238), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 key_mem_reg_2__120_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1144]), 
	.D(FE_PHN4819_n1148), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_2__88_ (.RN(FE_OFN45_reset_n), 
	.Q(key_mem[1112]), 
	.D(FE_PHN4915_n1180), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 key_mem_reg_2__56_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1080]), 
	.D(FE_PHN4667_n1212), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_2__24_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1048]), 
	.D(FE_PHN739_n1244), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_2__127_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1151]), 
	.D(FE_PHN4908_n1141), 
	.CK(clk_48Mhz__L6_N42));
   DFFRHQX1 key_mem_reg_2__95_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1119]), 
	.D(FE_PHN4934_n1173), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 key_mem_reg_2__63_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1087]), 
	.D(FE_PHN789_n1205), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 key_mem_reg_2__31_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1055]), 
	.D(FE_PHN4790_n1237), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 prev_key1_reg_reg_87_ (.Q(prev_key1_reg[87]), 
	.D(FE_PHN4990_n2333), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 prev_key1_reg_reg_86_ (.Q(prev_key1_reg[86]), 
	.D(FE_PHN4995_n2334), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 prev_key1_reg_reg_85_ (.Q(prev_key1_reg[85]), 
	.D(FE_PHN5016_n2335), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 prev_key1_reg_reg_84_ (.Q(prev_key1_reg[84]), 
	.D(FE_PHN5011_n2336), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 prev_key1_reg_reg_83_ (.Q(prev_key1_reg[83]), 
	.D(FE_PHN4989_n2337), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 prev_key1_reg_reg_82_ (.Q(prev_key1_reg[82]), 
	.D(FE_PHN4999_n2338), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 prev_key1_reg_reg_81_ (.Q(prev_key1_reg[81]), 
	.D(FE_PHN5004_n2339), 
	.CK(clk_48Mhz__L6_N11));
   DFFHQX1 prev_key1_reg_reg_80_ (.Q(prev_key1_reg[80]), 
	.D(FE_PHN5003_n2340), 
	.CK(clk_48Mhz__L6_N11));
   DFFHQX1 prev_key1_reg_reg_79_ (.Q(prev_key1_reg[79]), 
	.D(FE_PHN5007_n2341), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 prev_key1_reg_reg_78_ (.Q(prev_key1_reg[78]), 
	.D(FE_PHN5001_n2342), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 prev_key1_reg_reg_77_ (.Q(prev_key1_reg[77]), 
	.D(FE_PHN5000_n2343), 
	.CK(clk_48Mhz__L6_N27));
   DFFHQX1 prev_key1_reg_reg_76_ (.Q(prev_key1_reg[76]), 
	.D(FE_PHN5024_n2344), 
	.CK(clk_48Mhz__L6_N27));
   DFFHQX1 prev_key1_reg_reg_75_ (.Q(prev_key1_reg[75]), 
	.D(FE_PHN5012_n2345), 
	.CK(clk_48Mhz__L6_N23));
   DFFHQX1 prev_key1_reg_reg_74_ (.Q(prev_key1_reg[74]), 
	.D(FE_PHN5013_n2346), 
	.CK(clk_48Mhz__L6_N14));
   DFFHQX1 prev_key1_reg_reg_73_ (.Q(prev_key1_reg[73]), 
	.D(FE_PHN5002_n2347), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 prev_key1_reg_reg_72_ (.Q(prev_key1_reg[72]), 
	.D(FE_PHN5008_n2348), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 prev_key1_reg_reg_71_ (.Q(prev_key1_reg[71]), 
	.D(FE_PHN5019_n2349), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 prev_key1_reg_reg_70_ (.Q(prev_key1_reg[70]), 
	.D(FE_PHN1035_n2350), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 prev_key1_reg_reg_69_ (.Q(prev_key1_reg[69]), 
	.D(FE_PHN5034_n2351), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 prev_key1_reg_reg_68_ (.Q(prev_key1_reg[68]), 
	.D(FE_PHN5029_n2352), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 prev_key1_reg_reg_67_ (.Q(prev_key1_reg[67]), 
	.D(FE_PHN5026_n2353), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 prev_key1_reg_reg_66_ (.Q(prev_key1_reg[66]), 
	.D(FE_PHN5025_n2354), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 prev_key1_reg_reg_65_ (.Q(prev_key1_reg[65]), 
	.D(FE_PHN4998_n2355), 
	.CK(clk));
   DFFHQX1 prev_key1_reg_reg_64_ (.Q(prev_key1_reg[64]), 
	.D(FE_PHN5022_n2356), 
	.CK(clk_48Mhz__L6_N34));
   DFFRHQX1 rcon_reg_reg_4_ (.RN(FE_OFN55_reset_n), 
	.Q(rcon_reg[4]), 
	.D(n2426), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 rcon_reg_reg_5_ (.RN(FE_OFN55_reset_n), 
	.Q(rcon_reg[5]), 
	.D(FE_PHN4980_n2425), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 rcon_reg_reg_1_ (.RN(FE_OFN55_reset_n), 
	.Q(rcon_reg[1]), 
	.D(n2429), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 rcon_reg_reg_6_ (.RN(FE_OFN55_reset_n), 
	.Q(rcon_reg[6]), 
	.D(FE_PHN4701_n2424), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 key_mem_reg_0__119_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1399]), 
	.D(FE_PHN2493_n893), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_0__118_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1398]), 
	.D(FE_PHN2634_n894), 
	.CK(clk_48Mhz__L6_N42));
   DFFRHQX1 key_mem_reg_0__117_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1397]), 
	.D(FE_PHN2417_n895), 
	.CK(clk_48Mhz__L6_N16));
   DFFRHQX1 key_mem_reg_0__116_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1396]), 
	.D(FE_PHN2675_n896), 
	.CK(clk_48Mhz__L6_N12));
   DFFRHQX1 key_mem_reg_0__115_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1395]), 
	.D(FE_PHN2503_n897), 
	.CK(clk_48Mhz__L6_N12));
   DFFRHQX1 key_mem_reg_0__114_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1394]), 
	.D(FE_PHN2507_n898), 
	.CK(clk_48Mhz__L6_N26));
   DFFRHQX1 key_mem_reg_0__113_ (.RN(FE_OFN39_reset_n), 
	.Q(key_mem[1393]), 
	.D(FE_PHN2702_n899), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 key_mem_reg_0__112_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1392]), 
	.D(FE_PHN2581_n900), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_0__111_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1391]), 
	.D(FE_PHN2440_n901), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 key_mem_reg_0__110_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1390]), 
	.D(FE_PHN4775_n902), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 key_mem_reg_0__109_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1389]), 
	.D(FE_PHN2630_n903), 
	.CK(clk_48Mhz__L6_N22));
   DFFRHQX1 key_mem_reg_0__108_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1388]), 
	.D(FE_PHN2487_n904), 
	.CK(clk_48Mhz__L6_N26));
   DFFRHQX1 key_mem_reg_0__107_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1387]), 
	.D(FE_PHN2545_n905), 
	.CK(clk_48Mhz__L6_N22));
   DFFRHQX1 key_mem_reg_0__106_ (.RN(FE_OFN55_reset_n), 
	.Q(key_mem[1386]), 
	.D(FE_PHN2411_n906), 
	.CK(clk_48Mhz__L6_N26));
   DFFRHQX1 key_mem_reg_0__105_ (.RN(FE_OFN39_reset_n), 
	.Q(key_mem[1385]), 
	.D(FE_PHN2641_n907), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 key_mem_reg_0__104_ (.RN(FE_OFN42_reset_n), 
	.Q(key_mem[1384]), 
	.D(FE_PHN1066_n908), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 key_mem_reg_0__103_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1383]), 
	.D(FE_PHN2551_n909), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 key_mem_reg_0__102_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1382]), 
	.D(FE_PHN2587_n910), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 key_mem_reg_0__101_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1381]), 
	.D(FE_PHN2609_n911), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 key_mem_reg_0__100_ (.RN(FE_OFN55_reset_n), 
	.Q(key_mem[1380]), 
	.D(FE_PHN2480_n912), 
	.CK(clk_48Mhz__L6_N26));
   DFFRHQX1 key_mem_reg_0__99_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1379]), 
	.D(FE_PHN4222_n913), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 key_mem_reg_0__98_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1378]), 
	.D(FE_PHN2657_n914), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 key_mem_reg_0__97_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1377]), 
	.D(FE_PHN2690_n915), 
	.CK(clk_48Mhz__L6_N34));
   DFFRHQX1 key_mem_reg_0__96_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1376]), 
	.D(FE_PHN2616_n916), 
	.CK(clk_48Mhz__L6_N25));
   DFFRHQX1 key_mem_reg_0__87_ (.RN(FE_OFN55_reset_n), 
	.Q(key_mem[1367]), 
	.D(FE_PHN2723_n925), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 key_mem_reg_0__86_ (.RN(FE_OFN43_reset_n), 
	.Q(key_mem[1366]), 
	.D(FE_PHN2754_n926), 
	.CK(clk_48Mhz__L6_N33));
   DFFRHQX1 key_mem_reg_0__85_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1365]), 
	.D(FE_PHN2629_n927), 
	.CK(clk_48Mhz__L6_N20));
   DFFRHQX1 key_mem_reg_0__84_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1364]), 
	.D(FE_PHN2713_n928), 
	.CK(clk_48Mhz__L6_N20));
   DFFRHQX1 key_mem_reg_0__83_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1363]), 
	.D(FE_PHN2684_n929), 
	.CK(clk_48Mhz__L6_N16));
   DFFRHQX1 key_mem_reg_0__82_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1362]), 
	.D(FE_PHN2589_n930), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 key_mem_reg_0__81_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1361]), 
	.D(FE_PHN2772_n931), 
	.CK(clk_48Mhz__L6_N7));
   DFFRHQX1 key_mem_reg_0__80_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1360]), 
	.D(FE_PHN2742_n932), 
	.CK(clk_48Mhz__L6_N7));
   DFFRHQX1 key_mem_reg_0__79_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1359]), 
	.D(FE_PHN2555_n933), 
	.CK(clk_48Mhz__L6_N3));
   DFFRHQX1 key_mem_reg_0__78_ (.RN(FE_OFN42_reset_n), 
	.Q(key_mem[1358]), 
	.D(FE_PHN2563_n934), 
	.CK(clk_48Mhz__L6_N1));
   DFFRHQX1 key_mem_reg_0__77_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1357]), 
	.D(FE_PHN2784_n935), 
	.CK(clk_48Mhz__L6_N7));
   DFFRHQX1 key_mem_reg_0__76_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1356]), 
	.D(FE_PHN2590_n936), 
	.CK(clk_48Mhz__L6_N7));
   DFFRHQX1 key_mem_reg_0__75_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1355]), 
	.D(FE_PHN2698_n937), 
	.CK(clk_48Mhz__L6_N25));
   DFFRHQX1 key_mem_reg_0__74_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1354]), 
	.D(FE_PHN2418_n938), 
	.CK(clk));
   DFFRHQX1 key_mem_reg_0__73_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1353]), 
	.D(FE_PHN2731_n939), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 key_mem_reg_0__72_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1352]), 
	.D(FE_PHN2652_n940), 
	.CK(clk_48Mhz__L6_N3));
   DFFRHQX1 key_mem_reg_0__71_ (.RN(FE_OFN42_reset_n), 
	.Q(key_mem[1351]), 
	.D(FE_PHN2517_n941), 
	.CK(clk_48Mhz__L6_N1));
   DFFRHQX1 key_mem_reg_0__70_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1350]), 
	.D(FE_PHN2740_n942), 
	.CK(clk_48Mhz__L6_N25));
   DFFRHQX1 key_mem_reg_0__69_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1349]), 
	.D(FE_PHN2565_n943), 
	.CK(clk_48Mhz__L6_N28));
   DFFRHQX1 key_mem_reg_0__68_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1348]), 
	.D(FE_PHN938_n944), 
	.CK(clk_48Mhz__L6_N28));
   DFFRHQX1 key_mem_reg_0__67_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1347]), 
	.D(FE_PHN2614_n945), 
	.CK(clk_48Mhz__L6_N32));
   DFFRHQX1 key_mem_reg_0__66_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1346]), 
	.D(FE_PHN930_n946), 
	.CK(clk_48Mhz__L6_N34));
   DFFRHQX1 key_mem_reg_0__65_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1345]), 
	.D(FE_PHN4302_n947), 
	.CK(clk_48Mhz__L6_N28));
   DFFRHQX1 key_mem_reg_0__64_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1344]), 
	.D(FE_PHN4589_n948), 
	.CK(clk_48Mhz__L6_N32));
   DFFRHQX1 key_mem_reg_0__55_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1335]), 
	.D(FE_PHN2790_n957), 
	.CK(clk_48Mhz__L6_N13));
   DFFRHQX1 key_mem_reg_0__54_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1334]), 
	.D(FE_PHN2767_n958), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_0__53_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1333]), 
	.D(FE_PHN2605_n959), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_0__52_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1332]), 
	.D(FE_PHN2721_n960), 
	.CK(clk_48Mhz__L6_N13));
   DFFRHQX1 key_mem_reg_0__51_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1331]), 
	.D(FE_PHN2599_n961), 
	.CK(clk_48Mhz__L6_N17));
   DFFRHQX1 key_mem_reg_0__50_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1330]), 
	.D(FE_PHN718_n962), 
	.CK(clk_48Mhz__L6_N13));
   DFFRHQX1 key_mem_reg_0__49_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1329]), 
	.D(FE_PHN2722_n963), 
	.CK(clk_48Mhz__L6_N24));
   DFFRHQX1 key_mem_reg_0__48_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1328]), 
	.D(FE_PHN2405_n964), 
	.CK(clk_48Mhz__L6_N24));
   DFFRHQX1 key_mem_reg_0__47_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1327]), 
	.D(FE_PHN2779_n965), 
	.CK(clk_48Mhz__L6_N31));
   DFFRHQX1 key_mem_reg_0__46_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1326]), 
	.D(FE_PHN2433_n966), 
	.CK(clk_48Mhz__L6_N24));
   DFFRHQX1 key_mem_reg_0__45_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1325]), 
	.D(FE_PHN2540_n967), 
	.CK(clk_48Mhz__L6_N33));
   DFFRHQX1 key_mem_reg_0__44_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1324]), 
	.D(FE_PHN727_n968), 
	.CK(clk_48Mhz__L6_N31));
   DFFRHQX1 key_mem_reg_0__43_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1323]), 
	.D(FE_PHN2434_n969), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_0__42_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1322]), 
	.D(FE_PHN2564_n970), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_0__41_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1321]), 
	.D(FE_PHN1321_n971), 
	.CK(clk_48Mhz__L6_N32));
   DFFRHQX1 key_mem_reg_0__40_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1320]), 
	.D(FE_PHN1318_n972), 
	.CK(clk_48Mhz__L6_N24));
   DFFRHQX1 key_mem_reg_0__39_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1319]), 
	.D(FE_PHN2778_n973), 
	.CK(clk_48Mhz__L6_N28));
   DFFRHQX1 key_mem_reg_0__38_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1318]), 
	.D(FE_PHN2770_n974), 
	.CK(clk_48Mhz__L6_N3));
   DFFRHQX1 key_mem_reg_0__37_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1317]), 
	.D(FE_PHN708_n975), 
	.CK(clk_48Mhz__L6_N25));
   DFFRHQX1 key_mem_reg_0__36_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1316]), 
	.D(FE_PHN2509_n976), 
	.CK(clk_48Mhz__L6_N25));
   DFFRHQX1 key_mem_reg_0__35_ (.RN(FE_OFN45_reset_n), 
	.Q(key_mem[1315]), 
	.D(FE_PHN2720_n977), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 key_mem_reg_0__34_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1314]), 
	.D(FE_PHN719_n978), 
	.CK(clk_48Mhz__L6_N34));
   DFFRHQX1 key_mem_reg_0__33_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1313]), 
	.D(FE_PHN2530_n979), 
	.CK(clk));
   DFFRHQX1 key_mem_reg_0__32_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1312]), 
	.D(FE_PHN2495_n980), 
	.CK(clk));
   DFFRHQX1 key_mem_reg_0__23_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1303]), 
	.D(FE_PHN2640_n989), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 key_mem_reg_0__22_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1302]), 
	.D(FE_PHN937_n990), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_0__21_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1301]), 
	.D(FE_PHN1077_n991), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_0__20_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1300]), 
	.D(FE_PHN2786_n992), 
	.CK(clk_48Mhz__L6_N42));
   DFFRHQX1 key_mem_reg_0__19_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1299]), 
	.D(FE_PHN2703_n993), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_0__18_ (.RN(FE_OFN39_reset_n), 
	.Q(key_mem[1298]), 
	.D(FE_PHN928_n994), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 key_mem_reg_0__17_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1297]), 
	.D(FE_PHN2692_n995), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 key_mem_reg_0__16_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1296]), 
	.D(FE_PHN2481_n996), 
	.CK(clk_48Mhz__L6_N42));
   DFFRHQX1 key_mem_reg_0__15_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1295]), 
	.D(FE_PHN2758_n997), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 key_mem_reg_0__14_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1294]), 
	.D(FE_PHN2660_n998), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_0__13_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1293]), 
	.D(FE_PHN2685_n999), 
	.CK(clk_48Mhz__L6_N22));
   DFFRHQX1 key_mem_reg_0__12_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1292]), 
	.D(FE_PHN2460_n1000), 
	.CK(clk_48Mhz__L6_N18));
   DFFRHQX1 key_mem_reg_0__11_ (.RN(FE_OFN39_reset_n), 
	.Q(key_mem[1291]), 
	.D(FE_PHN2712_n1001), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 key_mem_reg_0__10_ (.RN(FE_OFN55_reset_n), 
	.Q(key_mem[1290]), 
	.D(FE_PHN2674_n1002), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 key_mem_reg_0__9_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1289]), 
	.D(FE_PHN2400_n1003), 
	.CK(clk));
   DFFRHQX1 key_mem_reg_0__8_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1288]), 
	.D(FE_PHN581_n1004), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 key_mem_reg_0__7_ (.RN(FE_OFN42_reset_n), 
	.Q(key_mem[1287]), 
	.D(FE_PHN2730_n1005), 
	.CK(clk_48Mhz__L6_N1));
   DFFRHQX1 key_mem_reg_0__6_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1286]), 
	.D(FE_PHN2459_n1006), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 key_mem_reg_0__5_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1285]), 
	.D(FE_PHN2687_n1007), 
	.CK(clk_48Mhz__L6_N13));
   DFFRHQX1 key_mem_reg_0__4_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1284]), 
	.D(FE_PHN2761_n1008), 
	.CK(clk_48Mhz__L6_N13));
   DFFRHQX1 key_mem_reg_0__3_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1283]), 
	.D(FE_PHN2759_n1009), 
	.CK(clk_48Mhz__L6_N31));
   DFFRHQX1 key_mem_reg_0__2_ (.RN(FE_OFN55_reset_n), 
	.Q(key_mem[1282]), 
	.D(FE_PHN2528_n1010), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 key_mem_reg_0__1_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1281]), 
	.D(FE_PHN2548_n1011), 
	.CK(clk_48Mhz__L6_N7));
   DFFRHQX1 key_mem_reg_0__0_ (.RN(FE_OFN42_reset_n), 
	.Q(key_mem[1280]), 
	.D(FE_PHN971_n1012), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 key_mem_reg_0__121_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1401]), 
	.D(FE_PHN950_n891), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 key_mem_reg_0__89_ (.RN(FE_OFN43_reset_n), 
	.Q(key_mem[1369]), 
	.D(FE_PHN628_n923), 
	.CK(clk_48Mhz__L6_N33));
   DFFRHQX1 key_mem_reg_0__57_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1337]), 
	.D(FE_PHN712_n955), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_0__25_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1305]), 
	.D(FE_PHN717_n987), 
	.CK(clk_48Mhz__L6_N18));
   DFFRHQX1 key_mem_reg_0__122_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1402]), 
	.D(FE_PHN2393_n890), 
	.CK(clk_48Mhz__L6_N22));
   DFFRHQX1 key_mem_reg_0__90_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1370]), 
	.D(FE_PHN2512_n922), 
	.CK(clk_48Mhz__L6_N16));
   DFFRHQX1 key_mem_reg_0__58_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1338]), 
	.D(FE_PHN2757_n954), 
	.CK(clk_48Mhz__L6_N17));
   DFFRHQX1 key_mem_reg_0__26_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1306]), 
	.D(FE_PHN2665_n986), 
	.CK(clk_48Mhz__L6_N19));
   DFFRHQX1 key_mem_reg_0__123_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1403]), 
	.D(FE_PHN2457_n889), 
	.CK(clk_48Mhz__L6_N19));
   DFFRHQX1 key_mem_reg_0__91_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1371]), 
	.D(FE_PHN2489_n921), 
	.CK(clk_48Mhz__L6_N16));
   DFFRHQX1 key_mem_reg_0__59_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1339]), 
	.D(FE_PHN731_n953), 
	.CK(clk_48Mhz__L6_N17));
   DFFRHQX1 key_mem_reg_0__27_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1307]), 
	.D(FE_PHN709_n985), 
	.CK(clk_48Mhz__L6_N19));
   DFFRHQX1 key_mem_reg_0__124_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1404]), 
	.D(FE_PHN994_n888), 
	.CK(clk_48Mhz__L6_N12));
   DFFRHQX1 key_mem_reg_0__92_ (.RN(FE_OFN43_reset_n), 
	.Q(key_mem[1372]), 
	.D(FE_PHN4751_n920), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 key_mem_reg_0__60_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1340]), 
	.D(FE_PHN2468_n952), 
	.CK(clk_48Mhz__L6_N33));
   DFFRHQX1 key_mem_reg_0__28_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1308]), 
	.D(FE_PHN2570_n984), 
	.CK(clk_48Mhz__L6_N22));
   DFFRHQX1 key_mem_reg_0__125_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1405]), 
	.D(FE_PHN2700_n887), 
	.CK(clk_48Mhz__L6_N12));
   DFFRHQX1 key_mem_reg_0__93_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1373]), 
	.D(FE_PHN2662_n919), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 key_mem_reg_0__61_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1341]), 
	.D(FE_PHN2475_n951), 
	.CK(clk_48Mhz__L6_N33));
   DFFRHQX1 key_mem_reg_0__29_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1309]), 
	.D(FE_PHN2602_n983), 
	.CK(clk_48Mhz__L6_N22));
   DFFRHQX1 key_mem_reg_0__126_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1406]), 
	.D(FE_PHN2777_n886), 
	.CK(clk_48Mhz__L6_N42));
   DFFRHQX1 key_mem_reg_0__94_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1374]), 
	.D(FE_PHN2788_n918), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 key_mem_reg_0__62_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1342]), 
	.D(FE_PHN2431_n950), 
	.CK(clk_48Mhz__L6_N32));
   DFFRHQX1 key_mem_reg_0__30_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1310]), 
	.D(FE_PHN2479_n982), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 key_mem_reg_0__120_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1400]), 
	.D(FE_PHN976_n892), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_0__88_ (.RN(FE_OFN45_reset_n), 
	.Q(key_mem[1368]), 
	.D(FE_PHN2465_n924), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 key_mem_reg_0__56_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1336]), 
	.D(FE_PHN2633_n956), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_0__24_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1304]), 
	.D(FE_PHN2556_n988), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_0__127_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1407]), 
	.D(FE_PHN2738_n885), 
	.CK(clk_48Mhz__L6_N42));
   DFFRHQX1 key_mem_reg_0__95_ (.RN(FE_OFN42_reset_n), 
	.Q(key_mem[1375]), 
	.D(FE_PHN631_n917), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 key_mem_reg_0__63_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1343]), 
	.D(FE_PHN2568_n949), 
	.CK(clk_48Mhz__L6_N32));
   DFFRHQX1 key_mem_reg_0__31_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1311]), 
	.D(FE_PHN4931_n981), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 key_mem_reg_1__119_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1271]), 
	.D(FE_PHN4873_n1021), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_1__118_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1270]), 
	.D(FE_PHN1096_n1022), 
	.CK(clk_48Mhz__L6_N42));
   DFFRHQX1 key_mem_reg_1__117_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1269]), 
	.D(FE_PHN1076_n1023), 
	.CK(clk_48Mhz__L6_N17));
   DFFRHQX1 key_mem_reg_1__116_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1268]), 
	.D(FE_PHN4204_n1024), 
	.CK(clk_48Mhz__L6_N16));
   DFFRHQX1 key_mem_reg_1__115_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1267]), 
	.D(FE_PHN4648_n1025), 
	.CK(clk_48Mhz__L6_N12));
   DFFRHQX1 key_mem_reg_1__114_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1266]), 
	.D(FE_PHN4619_n1026), 
	.CK(clk_48Mhz__L6_N16));
   DFFRHQX1 key_mem_reg_1__113_ (.RN(FE_OFN39_reset_n), 
	.Q(key_mem[1265]), 
	.D(FE_PHN4978_n1027), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 key_mem_reg_1__112_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1264]), 
	.D(FE_PHN4366_n1028), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_1__111_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1263]), 
	.D(FE_PHN1324_n1029), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 key_mem_reg_1__110_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1262]), 
	.D(FE_PHN1322_n1030), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_1__109_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1261]), 
	.D(FE_PHN4470_n1031), 
	.CK(clk_48Mhz__L6_N19));
   DFFRHQX1 key_mem_reg_1__108_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1260]), 
	.D(FE_PHN4191_n1032), 
	.CK(clk_48Mhz__L6_N26));
   DFFRHQX1 key_mem_reg_1__107_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1259]), 
	.D(FE_PHN4959_n1033), 
	.CK(clk_48Mhz__L6_N22));
   DFFRHQX1 key_mem_reg_1__106_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1258]), 
	.D(FE_PHN4538_n1034), 
	.CK(clk_48Mhz__L6_N26));
   DFFRHQX1 key_mem_reg_1__105_ (.RN(FE_OFN39_reset_n), 
	.Q(key_mem[1257]), 
	.D(FE_PHN4523_n1035), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 key_mem_reg_1__104_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1256]), 
	.D(FE_PHN4647_n1036), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 key_mem_reg_1__103_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1255]), 
	.D(FE_PHN4898_n1037), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 key_mem_reg_1__102_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1254]), 
	.D(FE_PHN4925_n1038), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 key_mem_reg_1__101_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1253]), 
	.D(FE_PHN4804_n1039), 
	.CK(clk_48Mhz__L6_N26));
   DFFRHQX1 key_mem_reg_1__100_ (.RN(FE_OFN55_reset_n), 
	.Q(key_mem[1252]), 
	.D(FE_PHN4226_n1040), 
	.CK(clk_48Mhz__L6_N26));
   DFFRHQX1 key_mem_reg_1__99_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1251]), 
	.D(FE_PHN1085_n1041), 
	.CK(clk_48Mhz__L6_N34));
   DFFRHQX1 key_mem_reg_1__98_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1250]), 
	.D(FE_PHN4287_n1042), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 key_mem_reg_1__97_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1249]), 
	.D(FE_PHN4778_n1043), 
	.CK(clk_48Mhz__L6_N34));
   DFFRHQX1 key_mem_reg_1__96_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1248]), 
	.D(FE_PHN4561_n1044), 
	.CK(clk_48Mhz__L6_N25));
   DFFRHQX1 key_mem_reg_1__87_ (.RN(FE_OFN55_reset_n), 
	.Q(key_mem[1239]), 
	.D(FE_PHN4789_n1053), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 key_mem_reg_1__86_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1238]), 
	.D(FE_PHN4234_n1054), 
	.CK(clk_48Mhz__L6_N33));
   DFFRHQX1 key_mem_reg_1__85_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1237]), 
	.D(FE_PHN970_n1055), 
	.CK(clk_48Mhz__L6_N20));
   DFFRHQX1 key_mem_reg_1__84_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1236]), 
	.D(FE_PHN4418_n1056), 
	.CK(clk_48Mhz__L6_N20));
   DFFRHQX1 key_mem_reg_1__83_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1235]), 
	.D(FE_PHN4539_n1057), 
	.CK(clk_48Mhz__L6_N16));
   DFFRHQX1 key_mem_reg_1__82_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1234]), 
	.D(FE_PHN4742_n1058), 
	.CK(clk_48Mhz__L6_N16));
   DFFRHQX1 key_mem_reg_1__81_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1233]), 
	.D(FE_PHN810_n1059), 
	.CK(clk));
   DFFRHQX1 key_mem_reg_1__80_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1232]), 
	.D(FE_PHN4328_n1060), 
	.CK(clk_48Mhz__L6_N7));
   DFFRHQX1 key_mem_reg_1__79_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1231]), 
	.D(FE_PHN4484_n1061), 
	.CK(clk_48Mhz__L6_N3));
   DFFRHQX1 key_mem_reg_1__78_ (.RN(FE_OFN42_reset_n), 
	.Q(key_mem[1230]), 
	.D(FE_PHN4958_n1062), 
	.CK(clk_48Mhz__L6_N1));
   DFFRHQX1 key_mem_reg_1__77_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1229]), 
	.D(FE_PHN4187_n1063), 
	.CK(clk_48Mhz__L6_N7));
   DFFRHQX1 key_mem_reg_1__76_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1228]), 
	.D(FE_PHN4413_n1064), 
	.CK(clk_48Mhz__L6_N7));
   DFFRHQX1 key_mem_reg_1__75_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1227]), 
	.D(FE_PHN4826_n1065), 
	.CK(clk_48Mhz__L6_N25));
   DFFRHQX1 key_mem_reg_1__74_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1226]), 
	.D(FE_PHN4800_n1066), 
	.CK(clk));
   DFFRHQX1 key_mem_reg_1__73_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1225]), 
	.D(FE_PHN4966_n1067), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 key_mem_reg_1__72_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1224]), 
	.D(FE_PHN4578_n1068), 
	.CK(clk_48Mhz__L6_N3));
   DFFRHQX1 key_mem_reg_1__71_ (.RN(FE_OFN42_reset_n), 
	.Q(key_mem[1223]), 
	.D(FE_PHN4653_n1069), 
	.CK(clk_48Mhz__L6_N1));
   DFFRHQX1 key_mem_reg_1__70_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1222]), 
	.D(FE_PHN4834_n1070), 
	.CK(clk_48Mhz__L6_N25));
   DFFRHQX1 key_mem_reg_1__69_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1221]), 
	.D(FE_PHN923_n1071), 
	.CK(clk_48Mhz__L6_N28));
   DFFRHQX1 key_mem_reg_1__68_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1220]), 
	.D(FE_PHN4627_n1072), 
	.CK(clk_48Mhz__L6_N28));
   DFFRHQX1 key_mem_reg_1__67_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1219]), 
	.D(FE_PHN4963_n1073), 
	.CK(clk_48Mhz__L6_N32));
   DFFRHQX1 key_mem_reg_1__66_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1218]), 
	.D(FE_PHN4296_n1074), 
	.CK(clk_48Mhz__L6_N34));
   DFFRHQX1 key_mem_reg_1__65_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1217]), 
	.D(FE_PHN2769_n1075), 
	.CK(clk_48Mhz__L6_N28));
   DFFRHQX1 key_mem_reg_1__64_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1216]), 
	.D(FE_PHN1011_n1076), 
	.CK(clk_48Mhz__L6_N34));
   DFFRHQX1 key_mem_reg_1__55_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1207]), 
	.D(FE_PHN4979_n1085), 
	.CK(clk_48Mhz__L6_N13));
   DFFRHQX1 key_mem_reg_1__54_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1206]), 
	.D(FE_PHN4889_n1086), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_1__53_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1205]), 
	.D(FE_PHN4860_n1087), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_1__52_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1204]), 
	.D(FE_PHN720_n1088), 
	.CK(clk_48Mhz__L6_N13));
   DFFRHQX1 key_mem_reg_1__51_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1203]), 
	.D(FE_PHN4471_n1089), 
	.CK(clk_48Mhz__L6_N17));
   DFFRHQX1 key_mem_reg_1__50_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1202]), 
	.D(FE_PHN4700_n1090), 
	.CK(clk_48Mhz__L6_N13));
   DFFRHQX1 key_mem_reg_1__49_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1201]), 
	.D(FE_PHN4822_n1091), 
	.CK(clk_48Mhz__L6_N24));
   DFFRHQX1 key_mem_reg_1__48_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1200]), 
	.D(FE_PHN4576_n1092), 
	.CK(clk_48Mhz__L6_N24));
   DFFRHQX1 key_mem_reg_1__47_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1199]), 
	.D(FE_PHN4740_n1093), 
	.CK(clk_48Mhz__L6_N31));
   DFFRHQX1 key_mem_reg_1__46_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1198]), 
	.D(FE_PHN4414_n1094), 
	.CK(clk_48Mhz__L6_N32));
   DFFRHQX1 key_mem_reg_1__45_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1197]), 
	.D(FE_PHN726_n1095), 
	.CK(clk_48Mhz__L6_N33));
   DFFRHQX1 key_mem_reg_1__44_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1196]), 
	.D(FE_PHN4311_n1096), 
	.CK(clk_48Mhz__L6_N31));
   DFFRHQX1 key_mem_reg_1__43_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1195]), 
	.D(FE_PHN4367_n1097), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_1__42_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1194]), 
	.D(FE_PHN4677_n1098), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_1__41_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1193]), 
	.D(FE_PHN4935_n1099), 
	.CK(clk_48Mhz__L6_N28));
   DFFRHQX1 key_mem_reg_1__40_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1192]), 
	.D(FE_PHN4831_n1100), 
	.CK(clk_48Mhz__L6_N24));
   DFFRHQX1 key_mem_reg_1__39_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1191]), 
	.D(FE_PHN4520_n1101), 
	.CK(clk_48Mhz__L6_N24));
   DFFRHQX1 key_mem_reg_1__38_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1190]), 
	.D(FE_PHN706_n1102), 
	.CK(clk_48Mhz__L6_N3));
   DFFRHQX1 key_mem_reg_1__37_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1189]), 
	.D(FE_PHN4777_n1103), 
	.CK(clk_48Mhz__L6_N25));
   DFFRHQX1 key_mem_reg_1__36_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1188]), 
	.D(FE_PHN4307_n1104), 
	.CK(clk_48Mhz__L6_N25));
   DFFRHQX1 key_mem_reg_1__35_ (.RN(FE_OFN45_reset_n), 
	.Q(key_mem[1187]), 
	.D(FE_PHN716_n1105), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 key_mem_reg_1__34_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1186]), 
	.D(FE_PHN4862_n1106), 
	.CK(clk_48Mhz__L6_N34));
   DFFRHQX1 key_mem_reg_1__33_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1185]), 
	.D(FE_PHN724_n1107), 
	.CK(clk));
   DFFRHQX1 key_mem_reg_1__32_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1184]), 
	.D(FE_PHN4649_n1108), 
	.CK(clk_48Mhz__L6_N7));
   DFFRHQX1 key_mem_reg_1__23_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1175]), 
	.D(FE_PHN4744_n1117), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 key_mem_reg_1__22_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1174]), 
	.D(FE_PHN4960_n1118), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_1__21_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1173]), 
	.D(FE_PHN4708_n1119), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_1__20_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1172]), 
	.D(FE_PHN4640_n1120), 
	.CK(clk_48Mhz__L6_N42));
   DFFRHQX1 key_mem_reg_1__19_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1171]), 
	.D(FE_PHN986_n1121), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_1__18_ (.RN(FE_OFN39_reset_n), 
	.Q(key_mem[1170]), 
	.D(FE_PHN4453_n1122), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 key_mem_reg_1__17_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1169]), 
	.D(FE_PHN4638_n1123), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 key_mem_reg_1__16_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1168]), 
	.D(FE_PHN963_n1124), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_1__15_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1167]), 
	.D(FE_PHN4694_n1125), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 key_mem_reg_1__14_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1166]), 
	.D(FE_PHN4932_n1126), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_1__13_ (.RN(FE_OFN39_reset_n), 
	.Q(key_mem[1165]), 
	.D(FE_PHN944_n1127), 
	.CK(clk_48Mhz__L6_N19));
   DFFRHQX1 key_mem_reg_1__12_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1164]), 
	.D(FE_PHN956_n1128), 
	.CK(clk_48Mhz__L6_N18));
   DFFRHQX1 key_mem_reg_1__11_ (.RN(FE_OFN39_reset_n), 
	.Q(key_mem[1163]), 
	.D(FE_PHN4769_n1129), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 key_mem_reg_1__10_ (.RN(FE_OFN55_reset_n), 
	.Q(key_mem[1162]), 
	.D(FE_PHN4680_n1130), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 key_mem_reg_1__9_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1161]), 
	.D(FE_PHN4710_n1131), 
	.CK(clk_48Mhz__L6_N7));
   DFFRHQX1 key_mem_reg_1__8_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1160]), 
	.D(FE_PHN586_n1132), 
	.CK(clk_48Mhz__L6_N34));
   DFFRHQX1 key_mem_reg_1__7_ (.RN(FE_OFN42_reset_n), 
	.Q(key_mem[1159]), 
	.D(FE_PHN4610_n1133), 
	.CK(clk_48Mhz__L6_N1));
   DFFRHQX1 key_mem_reg_1__6_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1158]), 
	.D(FE_PHN4841_n1134), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 key_mem_reg_1__5_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1157]), 
	.D(FE_PHN4528_n1135), 
	.CK(clk_48Mhz__L6_N17));
   DFFRHQX1 key_mem_reg_1__4_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1156]), 
	.D(FE_PHN4604_n1136), 
	.CK(clk_48Mhz__L6_N13));
   DFFRHQX1 key_mem_reg_1__3_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1155]), 
	.D(FE_PHN4904_n1137), 
	.CK(clk_48Mhz__L6_N31));
   DFFRHQX1 key_mem_reg_1__2_ (.RN(FE_OFN39_reset_n), 
	.Q(key_mem[1154]), 
	.D(FE_PHN4725_n1138), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 key_mem_reg_1__1_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1153]), 
	.D(FE_PHN4890_n1139), 
	.CK(clk_48Mhz__L6_N7));
   DFFRHQX1 key_mem_reg_1__0_ (.RN(FE_OFN42_reset_n), 
	.Q(key_mem[1152]), 
	.D(FE_PHN4400_n1140), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 key_mem_reg_1__121_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1273]), 
	.D(FE_PHN4752_n1019), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 key_mem_reg_1__89_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1241]), 
	.D(FE_PHN4403_n1051), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 key_mem_reg_1__57_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1209]), 
	.D(FE_PHN4460_n1083), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_1__25_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1177]), 
	.D(FE_PHN4846_n1115), 
	.CK(clk_48Mhz__L6_N18));
   DFFRHQX1 key_mem_reg_1__122_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1274]), 
	.D(FE_PHN4579_n1018), 
	.CK(clk_48Mhz__L6_N22));
   DFFRHQX1 key_mem_reg_1__90_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1242]), 
	.D(FE_PHN4540_n1050), 
	.CK(clk_48Mhz__L6_N16));
   DFFRHQX1 key_mem_reg_1__58_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1210]), 
	.D(FE_PHN589_n1082), 
	.CK(clk_48Mhz__L6_N17));
   DFFRHQX1 key_mem_reg_1__26_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1178]), 
	.D(FE_PHN713_n1114), 
	.CK(clk_48Mhz__L6_N19));
   DFFRHQX1 key_mem_reg_1__123_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1275]), 
	.D(FE_PHN982_n1017), 
	.CK(clk_48Mhz__L6_N19));
   DFFRHQX1 key_mem_reg_1__91_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1243]), 
	.D(FE_PHN4522_n1049), 
	.CK(clk_48Mhz__L6_N26));
   DFFRHQX1 key_mem_reg_1__59_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1211]), 
	.D(FE_PHN4252_n1081), 
	.CK(clk_48Mhz__L6_N17));
   DFFRHQX1 key_mem_reg_1__27_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1179]), 
	.D(FE_PHN4553_n1113), 
	.CK(clk_48Mhz__L6_N18));
   DFFRHQX1 key_mem_reg_1__124_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1276]), 
	.D(FE_PHN4357_n1016), 
	.CK(clk_48Mhz__L6_N12));
   DFFRHQX1 key_mem_reg_1__92_ (.RN(FE_OFN43_reset_n), 
	.Q(key_mem[1244]), 
	.D(FE_PHN638_n1048), 
	.CK(clk_48Mhz__L6_N33));
   DFFRHQX1 key_mem_reg_1__60_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1212]), 
	.D(FE_PHN4546_n1080), 
	.CK(clk_48Mhz__L6_N32));
   DFFRHQX1 key_mem_reg_1__28_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1180]), 
	.D(FE_PHN730_n1112), 
	.CK(clk_48Mhz__L6_N22));
   DFFRHQX1 key_mem_reg_1__125_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1277]), 
	.D(FE_PHN4573_n1015), 
	.CK(clk_48Mhz__L6_N12));
   DFFRHQX1 key_mem_reg_1__93_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1245]), 
	.D(FE_PHN4447_n1047), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 key_mem_reg_1__61_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1213]), 
	.D(FE_PHN4320_n1079), 
	.CK(clk_48Mhz__L6_N33));
   DFFRHQX1 key_mem_reg_1__29_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1181]), 
	.D(FE_PHN721_n1111), 
	.CK(clk_48Mhz__L6_N22));
   DFFRHQX1 key_mem_reg_1__126_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1278]), 
	.D(FE_PHN4465_n1014), 
	.CK(clk_48Mhz__L6_N42));
   DFFRHQX1 key_mem_reg_1__94_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1246]), 
	.D(FE_PHN4495_n1046), 
	.CK(clk_48Mhz__L6_N3));
   DFFRHQX1 key_mem_reg_1__62_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1214]), 
	.D(FE_PHN4770_n1078), 
	.CK(clk_48Mhz__L6_N32));
   DFFRHQX1 key_mem_reg_1__30_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1182]), 
	.D(FE_PHN4717_n1110), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 key_mem_reg_1__120_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1272]), 
	.D(FE_PHN4971_n1020), 
	.CK(clk_48Mhz__L6_N18));
   DFFRHQX1 key_mem_reg_1__88_ (.RN(FE_OFN45_reset_n), 
	.Q(key_mem[1240]), 
	.D(FE_PHN4983_n1052), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 key_mem_reg_1__56_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1208]), 
	.D(FE_PHN4501_n1084), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_1__24_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1176]), 
	.D(FE_PHN4969_n1116), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_1__127_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1279]), 
	.D(FE_PHN1084_n1013), 
	.CK(clk_48Mhz__L6_N42));
   DFFRHQX1 key_mem_reg_1__95_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1247]), 
	.D(FE_PHN4870_n1045), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 key_mem_reg_1__63_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1215]), 
	.D(FE_PHN4368_n1077), 
	.CK(clk_48Mhz__L6_N32));
   DFFRHQX1 key_mem_reg_1__31_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1183]), 
	.D(FE_PHN2696_n1109), 
	.CK(clk_48Mhz__L6_N42));
   DFFRHQX1 rcon_reg_reg_7_ (.RN(FE_OFN55_reset_n), 
	.Q(rcon_reg[7]), 
	.D(FE_PHN5047_n2431), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 ready_reg_reg (.RN(FE_OFN39_reset_n), 
	.Q(ready), 
	.D(FE_PHN1032_n2868), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 rcon_reg_reg_2_ (.RN(FE_OFN55_reset_n), 
	.Q(rcon_reg[2]), 
	.D(FE_PHN4895_n2428), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 rcon_reg_reg_3_ (.RN(FE_OFN55_reset_n), 
	.Q(rcon_reg[3]), 
	.D(FE_PHN3403_n2427), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 rcon_reg_reg_0_ (.RN(FE_OFN55_reset_n), 
	.Q(rcon_reg[0]), 
	.D(FE_PHN5073_n2430), 
	.CK(clk_48Mhz__L6_N21));
   DFFHQX1 key_mem_reg_6__119_ (.Q(key_mem[631]), 
	.D(FE_PHN2062_n1661), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_6__118_ (.Q(key_mem[630]), 
	.D(FE_PHN2268_n1662), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_6__117_ (.Q(key_mem[629]), 
	.D(FE_PHN2612_n1663), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_6__116_ (.Q(key_mem[628]), 
	.D(FE_PHN2291_n1664), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_6__115_ (.Q(key_mem[627]), 
	.D(FE_PHN2259_n1665), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_6__114_ (.Q(key_mem[626]), 
	.D(FE_PHN2106_n1666), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_6__113_ (.Q(key_mem[625]), 
	.D(FE_PHN1487_n1667), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_6__108_ (.Q(key_mem[620]), 
	.D(FE_PHN2295_n1672), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_6__107_ (.Q(key_mem[619]), 
	.D(FE_PHN2430_n1673), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_6__105_ (.Q(key_mem[617]), 
	.D(FE_PHN1643_n1675), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_6__103_ (.Q(key_mem[615]), 
	.D(FE_PHN2313_n1677), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_6__102_ (.Q(key_mem[614]), 
	.D(FE_PHN2073_n1678), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_6__101_ (.Q(key_mem[613]), 
	.D(FE_PHN2198_n1679), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 key_mem_reg_6__100_ (.Q(key_mem[612]), 
	.D(FE_PHN2454_n1680), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_6__99_ (.Q(key_mem[611]), 
	.D(FE_PHN2442_n1681), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_6__81_ (.Q(key_mem[593]), 
	.D(FE_PHN2270_n1682), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_6__76_ (.Q(key_mem[588]), 
	.D(FE_PHN2050_n1687), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_6__75_ (.Q(key_mem[587]), 
	.D(FE_PHN964_n1688), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_6__73_ (.Q(key_mem[585]), 
	.D(FE_PHN2116_n1690), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_6__71_ (.Q(key_mem[583]), 
	.D(FE_PHN2120_n1692), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_6__70_ (.Q(key_mem[582]), 
	.D(FE_PHN2255_n1693), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_6__69_ (.Q(key_mem[581]), 
	.D(FE_PHN2370_n1694), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_6__68_ (.Q(key_mem[580]), 
	.D(FE_PHN2529_n1695), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_6__67_ (.Q(key_mem[579]), 
	.D(FE_PHN2213_n1696), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_6__66_ (.Q(key_mem[578]), 
	.D(FE_PHN2426_n1697), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_6__65_ (.Q(key_mem[577]), 
	.D(FE_PHN2448_n1698), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_6__55_ (.Q(key_mem[567]), 
	.D(FE_PHN2541_n1708), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_6__54_ (.Q(key_mem[566]), 
	.D(FE_PHN2385_n1709), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_6__53_ (.Q(key_mem[565]), 
	.D(FE_PHN2081_n1710), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_6__52_ (.Q(key_mem[564]), 
	.D(FE_PHN2383_n1711), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_6__51_ (.Q(key_mem[563]), 
	.D(FE_PHN2063_n1712), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_6__50_ (.Q(key_mem[562]), 
	.D(FE_PHN2102_n1713), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_6__49_ (.Q(key_mem[561]), 
	.D(FE_PHN2156_n1714), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_6__44_ (.Q(key_mem[556]), 
	.D(FE_PHN2348_n1719), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_6__43_ (.Q(key_mem[555]), 
	.D(FE_PHN2238_n1720), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_6__41_ (.Q(key_mem[553]), 
	.D(FE_PHN2175_n1722), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_6__39_ (.Q(key_mem[551]), 
	.D(FE_PHN2153_n1724), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_6__38_ (.Q(key_mem[550]), 
	.D(FE_PHN2484_n1725), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_6__37_ (.Q(key_mem[549]), 
	.D(FE_PHN2331_n1726), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_6__36_ (.Q(key_mem[548]), 
	.D(FE_PHN2235_n1727), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_6__35_ (.Q(key_mem[547]), 
	.D(FE_PHN2306_n1728), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 key_mem_reg_6__34_ (.Q(key_mem[546]), 
	.D(FE_PHN2197_n1729), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_6__33_ (.Q(key_mem[545]), 
	.D(FE_PHN2582_n1730), 
	.CK(clk));
   DFFHQX1 key_mem_reg_6__23_ (.Q(key_mem[535]), 
	.D(FE_PHN2515_n1740), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_6__22_ (.Q(key_mem[534]), 
	.D(FE_PHN2365_n1741), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_6__21_ (.Q(key_mem[533]), 
	.D(FE_PHN2360_n1742), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_6__20_ (.Q(key_mem[532]), 
	.D(FE_PHN2402_n1743), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_6__19_ (.Q(key_mem[531]), 
	.D(FE_PHN4587_n1744), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_6__18_ (.Q(key_mem[530]), 
	.D(FE_PHN1640_n1745), 
	.CK(clk_48Mhz__L6_N46));
   DFFHQX1 key_mem_reg_6__17_ (.Q(key_mem[529]), 
	.D(FE_PHN2664_n1746), 
	.CK(clk_48Mhz__L6_N47));
   DFFHQX1 key_mem_reg_6__12_ (.Q(key_mem[524]), 
	.D(FE_PHN1732_n1751), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_6__11_ (.Q(key_mem[523]), 
	.D(FE_PHN1486_n1752), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_6__9_ (.Q(key_mem[521]), 
	.D(FE_PHN2219_n1754), 
	.CK(clk));
   DFFHQX1 key_mem_reg_6__7_ (.Q(key_mem[519]), 
	.D(FE_PHN2252_n1756), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_6__6_ (.Q(key_mem[518]), 
	.D(FE_PHN2311_n1757), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 key_mem_reg_6__5_ (.Q(key_mem[517]), 
	.D(FE_PHN4379_n1758), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_6__4_ (.Q(key_mem[516]), 
	.D(FE_PHN2166_n1759), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_6__3_ (.Q(key_mem[515]), 
	.D(FE_PHN2183_n1760), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_6__2_ (.Q(key_mem[514]), 
	.D(FE_PHN2516_n1761), 
	.CK(clk_48Mhz__L6_N14));
   DFFHQX1 key_mem_reg_6__1_ (.Q(key_mem[513]), 
	.D(FE_PHN2075_n1762), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_6__98_ (.Q(key_mem[610]), 
	.D(FE_PHN2056_n1764), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 key_mem_reg_6__97_ (.Q(key_mem[609]), 
	.D(FE_PHN2669_n1765), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_6__87_ (.Q(key_mem[599]), 
	.D(FE_PHN2637_n1775), 
	.CK(clk_48Mhz__L6_N21));
   DFFHQX1 key_mem_reg_6__86_ (.Q(key_mem[598]), 
	.D(FE_PHN2505_n1776), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_6__85_ (.Q(key_mem[597]), 
	.D(FE_PHN2335_n1777), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_6__84_ (.Q(key_mem[596]), 
	.D(FE_PHN2330_n1778), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_6__83_ (.Q(key_mem[595]), 
	.D(FE_PHN2249_n1779), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_6__82_ (.Q(key_mem[594]), 
	.D(FE_PHN2432_n1780), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_9__119_ (.Q(key_mem[247]), 
	.D(FE_PHN2668_n2045), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_9__118_ (.Q(key_mem[246]), 
	.D(FE_PHN4542_n2046), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_9__117_ (.Q(key_mem[245]), 
	.D(FE_PHN1768_n2047), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_9__116_ (.Q(key_mem[244]), 
	.D(FE_PHN1513_n2048), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_9__115_ (.Q(key_mem[243]), 
	.D(FE_PHN2526_n2049), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_9__114_ (.Q(key_mem[242]), 
	.D(FE_PHN1470_n2050), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_9__113_ (.Q(key_mem[241]), 
	.D(FE_PHN2427_n2051), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_9__108_ (.Q(key_mem[236]), 
	.D(FE_PHN1471_n2056), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_9__107_ (.Q(key_mem[235]), 
	.D(FE_PHN1567_n2057), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_9__105_ (.Q(key_mem[233]), 
	.D(FE_PHN2199_n2059), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_9__103_ (.Q(key_mem[231]), 
	.D(FE_PHN1046_n2061), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 key_mem_reg_9__102_ (.Q(key_mem[230]), 
	.D(FE_PHN2101_n2062), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_9__101_ (.Q(key_mem[229]), 
	.D(FE_PHN1485_n2063), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 key_mem_reg_9__100_ (.Q(key_mem[228]), 
	.D(FE_PHN1591_n2064), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_9__99_ (.Q(key_mem[227]), 
	.D(FE_PHN2600_n2065), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_9__69_ (.Q(key_mem[197]), 
	.D(FE_PHN2547_n2066), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_9__68_ (.Q(key_mem[196]), 
	.D(FE_PHN2251_n2067), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_9__67_ (.Q(key_mem[195]), 
	.D(FE_PHN2108_n2068), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_9__66_ (.Q(key_mem[194]), 
	.D(FE_PHN2042_n2069), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_9__65_ (.Q(key_mem[193]), 
	.D(FE_PHN2162_n2070), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_9__55_ (.Q(key_mem[183]), 
	.D(FE_PHN2359_n2080), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_9__54_ (.Q(key_mem[182]), 
	.D(FE_PHN2127_n2081), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_9__53_ (.Q(key_mem[181]), 
	.D(FE_PHN2202_n2082), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_9__52_ (.Q(key_mem[180]), 
	.D(FE_PHN2247_n2083), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_9__51_ (.Q(key_mem[179]), 
	.D(FE_PHN2553_n2084), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_9__50_ (.Q(key_mem[178]), 
	.D(FE_PHN2377_n2085), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_9__49_ (.Q(key_mem[177]), 
	.D(FE_PHN2308_n2086), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_9__44_ (.Q(key_mem[172]), 
	.D(FE_PHN4928_n2091), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_9__43_ (.Q(key_mem[171]), 
	.D(FE_PHN2040_n2092), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_9__41_ (.Q(key_mem[169]), 
	.D(FE_PHN2561_n2094), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_9__39_ (.Q(key_mem[167]), 
	.D(FE_PHN2155_n2096), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_9__38_ (.Q(key_mem[166]), 
	.D(FE_PHN2244_n2097), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_9__37_ (.Q(key_mem[165]), 
	.D(FE_PHN2041_n2098), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_9__36_ (.Q(key_mem[164]), 
	.D(FE_PHN2157_n2099), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_9__35_ (.Q(key_mem[163]), 
	.D(FE_PHN2254_n2100), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 key_mem_reg_9__34_ (.Q(key_mem[162]), 
	.D(FE_PHN2280_n2101), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_9__33_ (.Q(key_mem[161]), 
	.D(FE_PHN2340_n2102), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_9__23_ (.Q(key_mem[151]), 
	.D(FE_PHN2339_n2112), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_9__22_ (.Q(key_mem[150]), 
	.D(FE_PHN2344_n2113), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_9__21_ (.Q(key_mem[149]), 
	.D(FE_PHN4749_n2114), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_9__20_ (.Q(key_mem[148]), 
	.D(FE_PHN2519_n2115), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_9__19_ (.Q(key_mem[147]), 
	.D(FE_PHN2677_n2116), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_9__18_ (.Q(key_mem[146]), 
	.D(FE_PHN2560_n2117), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_9__17_ (.Q(key_mem[145]), 
	.D(FE_PHN2470_n2118), 
	.CK(clk_48Mhz__L6_N47));
   DFFHQX1 key_mem_reg_9__12_ (.Q(key_mem[140]), 
	.D(FE_PHN2506_n2123), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_9__11_ (.Q(key_mem[139]), 
	.D(FE_PHN1466_n2124), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_9__9_ (.Q(key_mem[137]), 
	.D(FE_PHN2227_n2126), 
	.CK(clk));
   DFFHQX1 key_mem_reg_9__7_ (.Q(key_mem[135]), 
	.D(FE_PHN2342_n2128), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_9__6_ (.Q(key_mem[134]), 
	.D(FE_PHN2204_n2129), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 key_mem_reg_9__5_ (.Q(key_mem[133]), 
	.D(FE_PHN2354_n2130), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_9__4_ (.Q(key_mem[132]), 
	.D(FE_PHN2248_n2131), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_9__3_ (.Q(key_mem[131]), 
	.D(FE_PHN2115_n2132), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_9__2_ (.Q(key_mem[130]), 
	.D(FE_PHN1617_n2133), 
	.CK(clk_48Mhz__L6_N21));
   DFFHQX1 key_mem_reg_9__1_ (.Q(key_mem[129]), 
	.D(FE_PHN2390_n2134), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_9__98_ (.Q(key_mem[226]), 
	.D(FE_PHN2180_n2136), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 key_mem_reg_9__97_ (.Q(key_mem[225]), 
	.D(FE_PHN2129_n2137), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_9__87_ (.Q(key_mem[215]), 
	.D(FE_PHN1509_n2147), 
	.CK(clk_48Mhz__L6_N21));
   DFFHQX1 key_mem_reg_9__86_ (.Q(key_mem[214]), 
	.D(FE_PHN2533_n2148), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_9__85_ (.Q(key_mem[213]), 
	.D(FE_PHN2728_n2149), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_9__84_ (.Q(key_mem[212]), 
	.D(FE_PHN2472_n2150), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_9__83_ (.Q(key_mem[211]), 
	.D(FE_PHN1629_n2151), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_9__82_ (.Q(key_mem[210]), 
	.D(FE_PHN2090_n2152), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_9__81_ (.Q(key_mem[209]), 
	.D(FE_PHN2392_n2153), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_9__76_ (.Q(key_mem[204]), 
	.D(FE_PHN2109_n2158), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_9__75_ (.Q(key_mem[203]), 
	.D(FE_PHN2424_n2159), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_9__73_ (.Q(key_mem[201]), 
	.D(FE_PHN2406_n2161), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_9__71_ (.Q(key_mem[199]), 
	.D(FE_PHN2152_n2163), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_9__70_ (.Q(key_mem[198]), 
	.D(FE_PHN2283_n2164), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_6__121_ (.Q(key_mem[633]), 
	.D(FE_PHN1534_n1659), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_9__121_ (.Q(key_mem[249]), 
	.D(FE_PHN2410_n2043), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_6__89_ (.Q(key_mem[601]), 
	.D(FE_PHN2181_n1773), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_9__89_ (.Q(key_mem[217]), 
	.D(FE_PHN2278_n2145), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_6__57_ (.Q(key_mem[569]), 
	.D(FE_PHN2089_n1706), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_9__57_ (.Q(key_mem[185]), 
	.D(FE_PHN2301_n2078), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_6__25_ (.Q(key_mem[537]), 
	.D(FE_PHN1510_n1738), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_9__25_ (.Q(key_mem[153]), 
	.D(FE_PHN2325_n2110), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_6__123_ (.Q(key_mem[635]), 
	.D(FE_PHN1592_n1657), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_9__123_ (.Q(key_mem[251]), 
	.D(FE_PHN2347_n2041), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_6__91_ (.Q(key_mem[603]), 
	.D(FE_PHN2054_n1771), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_9__91_ (.Q(key_mem[219]), 
	.D(FE_PHN1705_n2143), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_6__59_ (.Q(key_mem[571]), 
	.D(FE_PHN2151_n1704), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_9__59_ (.Q(key_mem[187]), 
	.D(FE_PHN1490_n2076), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_6__27_ (.Q(key_mem[539]), 
	.D(FE_PHN1246_n1736), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_9__27_ (.Q(key_mem[155]), 
	.D(FE_PHN2443_n2108), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_6__124_ (.Q(key_mem[636]), 
	.D(FE_PHN2142_n1656), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_9__124_ (.Q(key_mem[252]), 
	.D(FE_PHN2537_n2040), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_6__92_ (.Q(key_mem[604]), 
	.D(FE_PHN2282_n1770), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_9__92_ (.Q(key_mem[220]), 
	.D(FE_PHN2145_n2142), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_6__60_ (.Q(key_mem[572]), 
	.D(FE_PHN2546_n1703), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_9__60_ (.Q(key_mem[188]), 
	.D(FE_PHN2372_n2075), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_6__28_ (.Q(key_mem[540]), 
	.D(FE_PHN2436_n1735), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_9__28_ (.Q(key_mem[156]), 
	.D(FE_PHN1499_n2107), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_7__108_ (.Q(key_mem[492]), 
	.D(FE_PHN2397_n1783), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_7__107_ (.Q(key_mem[491]), 
	.D(FE_PHN2642_n1784), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_7__105_ (.Q(key_mem[489]), 
	.D(FE_PHN2008_n1786), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_7__103_ (.Q(key_mem[487]), 
	.D(FE_PHN2233_n1788), 
	.CK(clk_48Mhz__L6_N6));
   DFFHQX1 key_mem_reg_7__102_ (.Q(key_mem[486]), 
	.D(FE_PHN2169_n1789), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_7__101_ (.Q(key_mem[485]), 
	.D(FE_PHN2695_n1790), 
	.CK(clk_48Mhz__L6_N14));
   DFFHQX1 key_mem_reg_7__100_ (.Q(key_mem[484]), 
	.D(FE_PHN2337_n1791), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_7__99_ (.Q(key_mem[483]), 
	.D(FE_PHN2240_n1792), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_7__119_ (.Q(key_mem[503]), 
	.D(FE_PHN2256_n1801), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_7__118_ (.Q(key_mem[502]), 
	.D(FE_PHN2143_n1802), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_7__117_ (.Q(key_mem[501]), 
	.D(FE_PHN2221_n1803), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_7__116_ (.Q(key_mem[500]), 
	.D(FE_PHN2192_n1804), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_7__115_ (.Q(key_mem[499]), 
	.D(FE_PHN2051_n1805), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_7__114_ (.Q(key_mem[498]), 
	.D(FE_PHN2451_n1806), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_7__113_ (.Q(key_mem[497]), 
	.D(FE_PHN1673_n1807), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_7__11_ (.Q(key_mem[395]), 
	.D(FE_PHN2661_n1810), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_7__9_ (.Q(key_mem[393]), 
	.D(FE_PHN2716_n1812), 
	.CK(clk));
   DFFHQX1 key_mem_reg_7__7_ (.Q(key_mem[391]), 
	.D(FE_PHN2096_n1814), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_7__6_ (.Q(key_mem[390]), 
	.D(FE_PHN2409_n1815), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_7__5_ (.Q(key_mem[389]), 
	.D(FE_PHN2601_n1816), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_7__4_ (.Q(key_mem[388]), 
	.D(FE_PHN2242_n1817), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_7__3_ (.Q(key_mem[387]), 
	.D(FE_PHN2111_n1818), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_7__2_ (.Q(key_mem[386]), 
	.D(FE_PHN2371_n1819), 
	.CK(clk_48Mhz__L6_N21));
   DFFHQX1 key_mem_reg_7__1_ (.Q(key_mem[385]), 
	.D(FE_PHN2185_n1820), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_7__98_ (.Q(key_mem[482]), 
	.D(FE_PHN2438_n1822), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 key_mem_reg_7__97_ (.Q(key_mem[481]), 
	.D(FE_PHN2266_n1823), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_7__87_ (.Q(key_mem[471]), 
	.D(FE_PHN2092_n1833), 
	.CK(clk_48Mhz__L6_N21));
   DFFHQX1 key_mem_reg_7__86_ (.Q(key_mem[470]), 
	.D(FE_PHN2196_n1834), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_7__85_ (.Q(key_mem[469]), 
	.D(FE_PHN2149_n1835), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_7__84_ (.Q(key_mem[468]), 
	.D(FE_PHN2676_n1836), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_7__83_ (.Q(key_mem[467]), 
	.D(FE_PHN2413_n1837), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_7__82_ (.Q(key_mem[466]), 
	.D(FE_PHN2550_n1838), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_7__81_ (.Q(key_mem[465]), 
	.D(FE_PHN2705_n1839), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_7__76_ (.Q(key_mem[460]), 
	.D(FE_PHN2212_n1844), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_7__75_ (.Q(key_mem[459]), 
	.D(FE_PHN2483_n1845), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_7__73_ (.Q(key_mem[457]), 
	.D(FE_PHN2174_n1847), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_7__71_ (.Q(key_mem[455]), 
	.D(FE_PHN2130_n1849), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_7__70_ (.Q(key_mem[454]), 
	.D(FE_PHN2160_n1850), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_7__69_ (.Q(key_mem[453]), 
	.D(FE_PHN2321_n1851), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_7__68_ (.Q(key_mem[452]), 
	.D(FE_PHN2105_n1852), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_7__67_ (.Q(key_mem[451]), 
	.D(FE_PHN2711_n1853), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_7__66_ (.Q(key_mem[450]), 
	.D(FE_PHN2309_n1854), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_7__65_ (.Q(key_mem[449]), 
	.D(FE_PHN2099_n1855), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_7__55_ (.Q(key_mem[439]), 
	.D(FE_PHN2394_n1865), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_7__54_ (.Q(key_mem[438]), 
	.D(FE_PHN2243_n1866), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_7__53_ (.Q(key_mem[437]), 
	.D(FE_PHN4774_n1867), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_7__52_ (.Q(key_mem[436]), 
	.D(FE_PHN2230_n1868), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_7__51_ (.Q(key_mem[435]), 
	.D(FE_PHN2414_n1869), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_7__50_ (.Q(key_mem[434]), 
	.D(FE_PHN2382_n1870), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_7__49_ (.Q(key_mem[433]), 
	.D(FE_PHN2203_n1871), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_7__44_ (.Q(key_mem[428]), 
	.D(FE_PHN2284_n1876), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_7__43_ (.Q(key_mem[427]), 
	.D(FE_PHN2229_n1877), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_7__41_ (.Q(key_mem[425]), 
	.D(FE_PHN2750_n1879), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_7__39_ (.Q(key_mem[423]), 
	.D(FE_PHN2375_n1881), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_7__38_ (.Q(key_mem[422]), 
	.D(FE_PHN2461_n1882), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_7__37_ (.Q(key_mem[421]), 
	.D(FE_PHN2343_n1883), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_7__36_ (.Q(key_mem[420]), 
	.D(FE_PHN2490_n1884), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_7__35_ (.Q(key_mem[419]), 
	.D(FE_PHN2049_n1885), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 key_mem_reg_7__34_ (.Q(key_mem[418]), 
	.D(FE_PHN2701_n1886), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_7__33_ (.Q(key_mem[417]), 
	.D(FE_PHN2163_n1887), 
	.CK(clk));
   DFFHQX1 key_mem_reg_7__23_ (.Q(key_mem[407]), 
	.D(FE_PHN2474_n1897), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_7__22_ (.Q(key_mem[406]), 
	.D(FE_PHN2218_n1898), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_7__21_ (.Q(key_mem[405]), 
	.D(FE_PHN2368_n1899), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_7__20_ (.Q(key_mem[404]), 
	.D(FE_PHN2522_n1900), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_7__19_ (.Q(key_mem[403]), 
	.D(FE_PHN2320_n1901), 
	.CK(clk_48Mhz__L6_N47));
   DFFHQX1 key_mem_reg_7__18_ (.Q(key_mem[402]), 
	.D(FE_PHN1480_n1902), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_7__17_ (.Q(key_mem[401]), 
	.D(FE_PHN2513_n1903), 
	.CK(clk_48Mhz__L6_N47));
   DFFHQX1 key_mem_reg_7__12_ (.Q(key_mem[396]), 
	.D(FE_PHN1610_n1908), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_4__119_ (.Q(key_mem[887]), 
	.D(FE_PHN2554_n1400), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_4__118_ (.Q(key_mem[886]), 
	.D(FE_PHN2446_n1401), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_4__117_ (.Q(key_mem[885]), 
	.D(FE_PHN2549_n1402), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_4__116_ (.Q(key_mem[884]), 
	.D(FE_PHN2606_n1403), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_4__115_ (.Q(key_mem[883]), 
	.D(FE_PHN2463_n1404), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_4__114_ (.Q(key_mem[882]), 
	.D(FE_PHN2085_n1405), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_4__113_ (.Q(key_mem[881]), 
	.D(FE_PHN2164_n1406), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_4__108_ (.Q(key_mem[876]), 
	.D(FE_PHN2323_n1411), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_4__107_ (.Q(key_mem[875]), 
	.D(FE_PHN2082_n1412), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_4__105_ (.Q(key_mem[873]), 
	.D(FE_PHN2485_n1414), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_4__103_ (.Q(key_mem[871]), 
	.D(FE_PHN2046_n1416), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 key_mem_reg_4__102_ (.Q(key_mem[870]), 
	.D(FE_PHN2104_n1417), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 key_mem_reg_4__101_ (.Q(key_mem[869]), 
	.D(FE_PHN1578_n1418), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_4__100_ (.Q(key_mem[868]), 
	.D(FE_PHN1540_n1419), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_4__99_ (.Q(key_mem[867]), 
	.D(FE_PHN2190_n1420), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 key_mem_reg_4__23_ (.Q(key_mem[791]), 
	.D(FE_PHN2095_n1426), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_4__22_ (.Q(key_mem[790]), 
	.D(FE_PHN2644_n1427), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_4__21_ (.Q(key_mem[789]), 
	.D(FE_PHN2577_n1428), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_4__20_ (.Q(key_mem[788]), 
	.D(FE_PHN2285_n1429), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_4__19_ (.Q(key_mem[787]), 
	.D(FE_PHN2659_n1430), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_4__18_ (.Q(key_mem[786]), 
	.D(FE_PHN2542_n1431), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_4__17_ (.Q(key_mem[785]), 
	.D(FE_PHN2682_n1432), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_4__12_ (.Q(key_mem[780]), 
	.D(FE_PHN2353_n1437), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_4__11_ (.Q(key_mem[779]), 
	.D(FE_PHN1686_n1438), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_4__9_ (.Q(key_mem[777]), 
	.D(FE_PHN2200_n1440), 
	.CK(clk));
   DFFHQX1 key_mem_reg_4__7_ (.Q(key_mem[775]), 
	.D(FE_PHN2131_n1442), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_4__6_ (.Q(key_mem[774]), 
	.D(FE_PHN2262_n1443), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 key_mem_reg_4__5_ (.Q(key_mem[773]), 
	.D(FE_PHN2206_n1444), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_4__4_ (.Q(key_mem[772]), 
	.D(FE_PHN2611_n1445), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_4__3_ (.Q(key_mem[771]), 
	.D(FE_PHN2170_n1446), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_4__2_ (.Q(key_mem[770]), 
	.D(FE_PHN1541_n1447), 
	.CK(clk_48Mhz__L6_N21));
   DFFHQX1 key_mem_reg_4__1_ (.Q(key_mem[769]), 
	.D(FE_PHN2407_n1448), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_4__98_ (.Q(key_mem[866]), 
	.D(FE_PHN2107_n1450), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 key_mem_reg_4__97_ (.Q(key_mem[865]), 
	.D(FE_PHN2228_n1451), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_4__87_ (.Q(key_mem[855]), 
	.D(FE_PHN1664_n1461), 
	.CK(clk_48Mhz__L6_N21));
   DFFHQX1 key_mem_reg_4__86_ (.Q(key_mem[854]), 
	.D(FE_PHN2281_n1462), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_4__85_ (.Q(key_mem[853]), 
	.D(FE_PHN2263_n1463), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_4__84_ (.Q(key_mem[852]), 
	.D(FE_PHN2627_n1464), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_4__83_ (.Q(key_mem[851]), 
	.D(FE_PHN2362_n1465), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_4__82_ (.Q(key_mem[850]), 
	.D(FE_PHN2378_n1466), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_4__81_ (.Q(key_mem[849]), 
	.D(FE_PHN2272_n1467), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_4__76_ (.Q(key_mem[844]), 
	.D(FE_PHN2391_n1472), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_4__75_ (.Q(key_mem[843]), 
	.D(FE_PHN2289_n1473), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_4__73_ (.Q(key_mem[841]), 
	.D(FE_PHN2312_n1475), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_4__71_ (.Q(key_mem[839]), 
	.D(FE_PHN2603_n1477), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_4__70_ (.Q(key_mem[838]), 
	.D(FE_PHN2492_n1478), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_4__69_ (.Q(key_mem[837]), 
	.D(FE_PHN2650_n1479), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_4__68_ (.Q(key_mem[836]), 
	.D(FE_PHN2305_n1480), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_4__67_ (.Q(key_mem[835]), 
	.D(FE_PHN3881_n1481), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_4__66_ (.Q(key_mem[834]), 
	.D(FE_PHN2191_n1482), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_4__65_ (.Q(key_mem[833]), 
	.D(FE_PHN2395_n1483), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_4__55_ (.Q(key_mem[823]), 
	.D(FE_PHN4514_n1493), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_4__54_ (.Q(key_mem[822]), 
	.D(FE_PHN2223_n1494), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_4__53_ (.Q(key_mem[821]), 
	.D(FE_PHN2525_n1495), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_4__52_ (.Q(key_mem[820]), 
	.D(FE_PHN2079_n1496), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_4__51_ (.Q(key_mem[819]), 
	.D(FE_PHN2179_n1497), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_4__50_ (.Q(key_mem[818]), 
	.D(FE_PHN2066_n1498), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_4__49_ (.Q(key_mem[817]), 
	.D(FE_PHN2080_n1499), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_4__44_ (.Q(key_mem[812]), 
	.D(FE_PHN2356_n1504), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_4__43_ (.Q(key_mem[811]), 
	.D(FE_PHN4327_n1505), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_4__41_ (.Q(key_mem[809]), 
	.D(FE_PHN2317_n1507), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_4__39_ (.Q(key_mem[807]), 
	.D(FE_PHN2237_n1509), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_4__38_ (.Q(key_mem[806]), 
	.D(FE_PHN4211_n1510), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_4__37_ (.Q(key_mem[805]), 
	.D(FE_PHN2039_n1511), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_4__36_ (.Q(key_mem[804]), 
	.D(FE_PHN2322_n1512), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_4__35_ (.Q(key_mem[803]), 
	.D(FE_PHN2404_n1513), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 key_mem_reg_4__34_ (.Q(key_mem[802]), 
	.D(FE_PHN2326_n1514), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_4__33_ (.Q(key_mem[801]), 
	.D(FE_PHN2562_n1515), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_10__119_ (.Q(key_mem[119]), 
	.D(FE_PHN2456_n2173), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_10__118_ (.Q(key_mem[118]), 
	.D(FE_PHN2504_n2174), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_10__117_ (.Q(key_mem[117]), 
	.D(FE_PHN2140_n2175), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_10__116_ (.Q(key_mem[116]), 
	.D(FE_PHN2576_n2176), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_10__115_ (.Q(key_mem[115]), 
	.D(FE_PHN2310_n2177), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_10__114_ (.Q(key_mem[114]), 
	.D(FE_PHN2211_n2178), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_10__113_ (.Q(key_mem[113]), 
	.D(FE_PHN1782_n2179), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_10__108_ (.Q(key_mem[108]), 
	.D(FE_PHN2408_n2184), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_10__107_ (.Q(key_mem[107]), 
	.D(FE_PHN1728_n2185), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_10__105_ (.Q(key_mem[105]), 
	.D(FE_PHN1548_n2187), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_10__103_ (.Q(key_mem[103]), 
	.D(FE_PHN4215_n2189), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_10__102_ (.Q(key_mem[102]), 
	.D(FE_PHN2168_n2190), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_10__101_ (.Q(key_mem[101]), 
	.D(FE_PHN2520_n2191), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 key_mem_reg_10__100_ (.Q(key_mem[100]), 
	.D(FE_PHN2253_n2192), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_10__99_ (.Q(key_mem[99]), 
	.D(FE_PHN2201_n2193), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 key_mem_reg_10__98_ (.Q(key_mem[98]), 
	.D(FE_PHN2387_n2194), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 key_mem_reg_10__97_ (.Q(key_mem[97]), 
	.D(FE_PHN2208_n2195), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_10__87_ (.Q(key_mem[87]), 
	.D(FE_PHN1665_n2205), 
	.CK(clk_48Mhz__L6_N21));
   DFFHQX1 key_mem_reg_10__86_ (.Q(key_mem[86]), 
	.D(FE_PHN2137_n2206), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_10__85_ (.Q(key_mem[85]), 
	.D(FE_PHN2439_n2207), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_10__84_ (.Q(key_mem[84]), 
	.D(FE_PHN2476_n2208), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_10__83_ (.Q(key_mem[83]), 
	.D(FE_PHN2471_n2209), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_10__82_ (.Q(key_mem[82]), 
	.D(FE_PHN2159_n2210), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_10__81_ (.Q(key_mem[81]), 
	.D(FE_PHN2070_n2211), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_10__76_ (.Q(key_mem[76]), 
	.D(FE_PHN2388_n2216), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_10__75_ (.Q(key_mem[75]), 
	.D(FE_PHN2333_n2217), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_10__73_ (.Q(key_mem[73]), 
	.D(FE_PHN2220_n2219), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_10__71_ (.Q(key_mem[71]), 
	.D(FE_PHN2052_n2221), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_10__70_ (.Q(key_mem[70]), 
	.D(FE_PHN2367_n2222), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_10__69_ (.Q(key_mem[69]), 
	.D(FE_PHN2626_n2223), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_10__68_ (.Q(key_mem[68]), 
	.D(FE_PHN2226_n2224), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_10__67_ (.Q(key_mem[67]), 
	.D(FE_PHN2329_n2225), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_10__66_ (.Q(key_mem[66]), 
	.D(FE_PHN2374_n2226), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_10__65_ (.Q(key_mem[65]), 
	.D(FE_PHN2352_n2227), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_10__55_ (.Q(key_mem[55]), 
	.D(FE_PHN2146_n2237), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_10__54_ (.Q(key_mem[54]), 
	.D(FE_PHN2292_n2238), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_10__53_ (.Q(key_mem[53]), 
	.D(FE_PHN2535_n2239), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_10__52_ (.Q(key_mem[52]), 
	.D(FE_PHN2258_n2240), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_10__51_ (.Q(key_mem[51]), 
	.D(FE_PHN2597_n2241), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_10__50_ (.Q(key_mem[50]), 
	.D(FE_PHN2184_n2242), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_10__49_ (.Q(key_mem[49]), 
	.D(FE_PHN2067_n2243), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_10__44_ (.Q(key_mem[44]), 
	.D(FE_PHN2502_n2248), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_10__43_ (.Q(key_mem[43]), 
	.D(FE_PHN2628_n2249), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_10__41_ (.Q(key_mem[41]), 
	.D(FE_PHN2114_n2251), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_10__39_ (.Q(key_mem[39]), 
	.D(FE_PHN2521_n2253), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_10__38_ (.Q(key_mem[38]), 
	.D(FE_PHN2524_n2254), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_10__37_ (.Q(key_mem[37]), 
	.D(FE_PHN2225_n2255), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_10__36_ (.Q(key_mem[36]), 
	.D(FE_PHN2195_n2256), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_10__35_ (.Q(key_mem[35]), 
	.D(FE_PHN2307_n2257), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 key_mem_reg_10__34_ (.Q(key_mem[34]), 
	.D(FE_PHN2488_n2258), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_10__33_ (.Q(key_mem[33]), 
	.D(FE_PHN2119_n2259), 
	.CK(clk));
   DFFHQX1 key_mem_reg_10__23_ (.Q(key_mem[23]), 
	.D(FE_PHN2386_n2269), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_10__22_ (.Q(key_mem[22]), 
	.D(FE_PHN2346_n2270), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_10__21_ (.Q(key_mem[21]), 
	.D(FE_PHN2579_n2271), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_10__20_ (.Q(key_mem[20]), 
	.D(FE_PHN2286_n2272), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_10__19_ (.Q(key_mem[19]), 
	.D(FE_PHN2139_n2273), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_10__18_ (.Q(key_mem[18]), 
	.D(FE_PHN2222_n2274), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_10__17_ (.Q(key_mem[17]), 
	.D(FE_PHN2455_n2275), 
	.CK(clk_48Mhz__L6_N47));
   DFFHQX1 key_mem_reg_10__12_ (.Q(key_mem[12]), 
	.D(FE_PHN1648_n2280), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_10__11_ (.Q(key_mem[11]), 
	.D(FE_PHN1526_n2281), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_10__9_ (.Q(key_mem[9]), 
	.D(FE_PHN2269_n2283), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_10__7_ (.Q(key_mem[7]), 
	.D(FE_PHN2194_n2285), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_10__6_ (.Q(key_mem[6]), 
	.D(FE_PHN2072_n2286), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 key_mem_reg_10__5_ (.Q(key_mem[5]), 
	.D(FE_PHN4184_n2287), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_10__4_ (.Q(key_mem[4]), 
	.D(FE_PHN2176_n2288), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_10__3_ (.Q(key_mem[3]), 
	.D(FE_PHN2573_n2289), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_10__2_ (.Q(key_mem[2]), 
	.D(FE_PHN2621_n2290), 
	.CK(clk_48Mhz__L6_N14));
   DFFHQX1 key_mem_reg_10__1_ (.Q(key_mem[1]), 
	.D(FE_PHN2552_n2291), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_4__121_ (.Q(key_mem[889]), 
	.D(FE_PHN2401_n1398), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_7__121_ (.Q(key_mem[505]), 
	.D(FE_PHN2009_n1799), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_10__121_ (.Q(key_mem[121]), 
	.D(FE_PHN1599_n2171), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_4__89_ (.Q(key_mem[857]), 
	.D(FE_PHN2059_n1459), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_7__89_ (.Q(key_mem[473]), 
	.D(FE_PHN2421_n1831), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_10__89_ (.Q(key_mem[89]), 
	.D(FE_PHN2345_n2203), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_4__57_ (.Q(key_mem[825]), 
	.D(FE_PHN2112_n1491), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_7__57_ (.Q(key_mem[441]), 
	.D(FE_PHN2214_n1863), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_10__57_ (.Q(key_mem[57]), 
	.D(FE_PHN2048_n2235), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_4__25_ (.Q(key_mem[793]), 
	.D(FE_PHN2358_n1523), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_7__25_ (.Q(key_mem[409]), 
	.D(FE_PHN1737_n1895), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_10__25_ (.Q(key_mem[25]), 
	.D(FE_PHN1837_n2267), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_4__123_ (.Q(key_mem[891]), 
	.D(FE_PHN2087_n1425), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_7__123_ (.Q(key_mem[507]), 
	.D(FE_PHN2435_n1797), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_10__123_ (.Q(key_mem[123]), 
	.D(FE_PHN1651_n2169), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_4__91_ (.Q(key_mem[859]), 
	.D(FE_PHN2349_n1457), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_7__91_ (.Q(key_mem[475]), 
	.D(FE_PHN2069_n1829), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_10__91_ (.Q(key_mem[91]), 
	.D(FE_PHN2260_n2201), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_4__59_ (.Q(key_mem[827]), 
	.D(FE_PHN2154_n1489), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_7__59_ (.Q(key_mem[443]), 
	.D(FE_PHN2498_n1861), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_10__59_ (.Q(key_mem[59]), 
	.D(FE_PHN2379_n2233), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_4__27_ (.Q(key_mem[795]), 
	.D(FE_PHN2265_n1521), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_7__27_ (.Q(key_mem[411]), 
	.D(FE_PHN2338_n1893), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_10__27_ (.Q(key_mem[27]), 
	.D(FE_PHN1558_n2265), 
	.CK(clk_48Mhz__L6_N19));
   DFFHQX1 key_mem_reg_4__124_ (.Q(key_mem[892]), 
	.D(FE_PHN2133_n1424), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_7__124_ (.Q(key_mem[508]), 
	.D(FE_PHN2065_n1796), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_10__124_ (.Q(key_mem[124]), 
	.D(FE_PHN2094_n2168), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_4__92_ (.Q(key_mem[860]), 
	.D(FE_PHN2224_n1456), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_7__92_ (.Q(key_mem[476]), 
	.D(FE_PHN2369_n1828), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_10__92_ (.Q(key_mem[92]), 
	.D(FE_PHN2177_n2200), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_4__60_ (.Q(key_mem[828]), 
	.D(FE_PHN2299_n1488), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_7__60_ (.Q(key_mem[444]), 
	.D(FE_PHN2315_n1860), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_10__60_ (.Q(key_mem[60]), 
	.D(FE_PHN2508_n2232), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_4__28_ (.Q(key_mem[796]), 
	.D(FE_PHN1647_n1520), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_7__28_ (.Q(key_mem[412]), 
	.D(FE_PHN2447_n1892), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_10__28_ (.Q(key_mem[28]), 
	.D(FE_PHN1566_n2264), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_8__119_ (.Q(key_mem[375]), 
	.D(FE_PHN4392_n1917), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_8__118_ (.Q(key_mem[374]), 
	.D(FE_PHN4586_n1918), 
	.CK(clk_48Mhz__L6_N43));
   DFFHQX1 key_mem_reg_8__117_ (.Q(key_mem[373]), 
	.D(FE_PHN4016_n1919), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_8__116_ (.Q(key_mem[372]), 
	.D(FE_PHN4083_n1920), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_8__115_ (.Q(key_mem[371]), 
	.D(FE_PHN3917_n1921), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_8__114_ (.Q(key_mem[370]), 
	.D(FE_PHN4786_n1922), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_8__113_ (.Q(key_mem[369]), 
	.D(FE_PHN4111_n1923), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_8__108_ (.Q(key_mem[364]), 
	.D(FE_PHN4042_n1928), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_8__107_ (.Q(key_mem[363]), 
	.D(FE_PHN4691_n1929), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_8__105_ (.Q(key_mem[361]), 
	.D(FE_PHN4271_n1931), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_8__103_ (.Q(key_mem[359]), 
	.D(FE_PHN4914_n1933), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 key_mem_reg_8__102_ (.Q(key_mem[358]), 
	.D(FE_PHN4594_n1934), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_8__101_ (.Q(key_mem[357]), 
	.D(FE_PHN4729_n1935), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_8__100_ (.Q(key_mem[356]), 
	.D(FE_PHN4505_n1936), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_8__99_ (.Q(key_mem[355]), 
	.D(FE_PHN4154_n1937), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_8__39_ (.Q(key_mem[295]), 
	.D(FE_PHN3846_n1939), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_8__38_ (.Q(key_mem[294]), 
	.D(FE_PHN4741_n1940), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_8__37_ (.Q(key_mem[293]), 
	.D(FE_PHN4059_n1941), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_8__36_ (.Q(key_mem[292]), 
	.D(FE_PHN4468_n1942), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_8__35_ (.Q(key_mem[291]), 
	.D(FE_PHN4866_n1943), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 key_mem_reg_8__34_ (.Q(key_mem[290]), 
	.D(FE_PHN4693_n1944), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_8__33_ (.Q(key_mem[289]), 
	.D(FE_PHN3786_n1945), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_8__23_ (.Q(key_mem[279]), 
	.D(FE_PHN4410_n1955), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_8__22_ (.Q(key_mem[278]), 
	.D(FE_PHN4388_n1956), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_8__21_ (.Q(key_mem[277]), 
	.D(FE_PHN3980_n1957), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_8__20_ (.Q(key_mem[276]), 
	.D(FE_PHN4168_n1958), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_8__19_ (.Q(key_mem[275]), 
	.D(FE_PHN4652_n1959), 
	.CK(clk_48Mhz__L6_N47));
   DFFHQX1 key_mem_reg_8__18_ (.Q(key_mem[274]), 
	.D(FE_PHN4411_n1960), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_8__17_ (.Q(key_mem[273]), 
	.D(FE_PHN4227_n1961), 
	.CK(clk_48Mhz__L6_N47));
   DFFHQX1 key_mem_reg_8__12_ (.Q(key_mem[268]), 
	.D(FE_PHN4563_n1966), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_8__11_ (.Q(key_mem[267]), 
	.D(FE_PHN1311_n1967), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_8__9_ (.Q(key_mem[265]), 
	.D(FE_PHN4437_n1969), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_8__7_ (.Q(key_mem[263]), 
	.D(FE_PHN4422_n1971), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_8__6_ (.Q(key_mem[262]), 
	.D(FE_PHN4601_n1972), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_8__5_ (.Q(key_mem[261]), 
	.D(FE_PHN4818_n1973), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_8__4_ (.Q(key_mem[260]), 
	.D(FE_PHN4491_n1974), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_8__3_ (.Q(key_mem[259]), 
	.D(FE_PHN4062_n1975), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_8__2_ (.Q(key_mem[258]), 
	.D(FE_PHN4869_n1976), 
	.CK(clk_48Mhz__L6_N14));
   DFFHQX1 key_mem_reg_8__1_ (.Q(key_mem[257]), 
	.D(FE_PHN4706_n1977), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_8__98_ (.Q(key_mem[354]), 
	.D(FE_PHN4745_n1979), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 key_mem_reg_8__97_ (.Q(key_mem[353]), 
	.D(FE_PHN4773_n1980), 
	.CK(clk));
   DFFHQX1 key_mem_reg_8__87_ (.Q(key_mem[343]), 
	.D(FE_PHN4722_n1990), 
	.CK(clk_48Mhz__L6_N21));
   DFFHQX1 key_mem_reg_8__86_ (.Q(key_mem[342]), 
	.D(FE_PHN4261_n1991), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_8__85_ (.Q(key_mem[341]), 
	.D(FE_PHN4675_n1992), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_8__84_ (.Q(key_mem[340]), 
	.D(FE_PHN4459_n1993), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_8__83_ (.Q(key_mem[339]), 
	.D(FE_PHN3646_n1994), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_8__82_ (.Q(key_mem[338]), 
	.D(FE_PHN4207_n1995), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_8__81_ (.Q(key_mem[337]), 
	.D(FE_PHN4210_n1996), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_8__76_ (.Q(key_mem[332]), 
	.D(FE_PHN3909_n2001), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_8__75_ (.Q(key_mem[331]), 
	.D(FE_PHN4066_n2002), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_8__73_ (.Q(key_mem[329]), 
	.D(FE_PHN4747_n2004), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_8__71_ (.Q(key_mem[327]), 
	.D(FE_PHN3961_n2006), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_8__70_ (.Q(key_mem[326]), 
	.D(FE_PHN4570_n2007), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_8__69_ (.Q(key_mem[325]), 
	.D(FE_PHN4346_n2008), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_8__68_ (.Q(key_mem[324]), 
	.D(FE_PHN4421_n2009), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_8__67_ (.Q(key_mem[323]), 
	.D(FE_PHN4562_n2010), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_8__66_ (.Q(key_mem[322]), 
	.D(FE_PHN4683_n2011), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_8__65_ (.Q(key_mem[321]), 
	.D(FE_PHN4248_n2012), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_8__55_ (.Q(key_mem[311]), 
	.D(FE_PHN4784_n2022), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_8__54_ (.Q(key_mem[310]), 
	.D(FE_PHN4329_n2023), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_8__53_ (.Q(key_mem[309]), 
	.D(FE_PHN4759_n2024), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_8__52_ (.Q(key_mem[308]), 
	.D(FE_PHN4322_n2025), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_8__51_ (.Q(key_mem[307]), 
	.D(FE_PHN4272_n2026), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_8__50_ (.Q(key_mem[306]), 
	.D(FE_PHN4292_n2027), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_8__49_ (.Q(key_mem[305]), 
	.D(FE_PHN4028_n2028), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_8__44_ (.Q(key_mem[300]), 
	.D(FE_PHN4728_n2033), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_8__43_ (.Q(key_mem[299]), 
	.D(FE_PHN3958_n2034), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_8__41_ (.Q(key_mem[297]), 
	.D(FE_PHN4835_n2036), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_5__119_ (.Q(key_mem[759]), 
	.D(FE_PHN4681_n1533), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_5__118_ (.Q(key_mem[758]), 
	.D(FE_PHN4548_n1534), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_5__117_ (.Q(key_mem[757]), 
	.D(FE_PHN4394_n1535), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_5__116_ (.Q(key_mem[756]), 
	.D(FE_PHN4486_n1536), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_5__115_ (.Q(key_mem[755]), 
	.D(FE_PHN4933_n1537), 
	.CK(clk_48Mhz__L6_N12));
   DFFHQX1 key_mem_reg_5__114_ (.Q(key_mem[754]), 
	.D(FE_PHN4633_n1538), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_5__113_ (.Q(key_mem[753]), 
	.D(FE_PHN1662_n1539), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_5__108_ (.Q(key_mem[748]), 
	.D(FE_PHN4035_n1544), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_5__107_ (.Q(key_mem[747]), 
	.D(FE_PHN1582_n1545), 
	.CK(clk_48Mhz__L6_N22));
   DFFHQX1 key_mem_reg_5__105_ (.Q(key_mem[745]), 
	.D(FE_PHN1733_n1547), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_5__103_ (.Q(key_mem[743]), 
	.D(FE_PHN3960_n1549), 
	.CK(clk_48Mhz__L6_N6));
   DFFHQX1 key_mem_reg_5__102_ (.Q(key_mem[742]), 
	.D(FE_PHN4791_n1550), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 key_mem_reg_5__101_ (.Q(key_mem[741]), 
	.D(FE_PHN4688_n1551), 
	.CK(clk_48Mhz__L6_N14));
   DFFHQX1 key_mem_reg_5__100_ (.Q(key_mem[740]), 
	.D(FE_PHN1681_n1552), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 key_mem_reg_5__99_ (.Q(key_mem[739]), 
	.D(FE_PHN4679_n1553), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_5__52_ (.Q(key_mem[692]), 
	.D(FE_PHN4399_n1554), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_5__51_ (.Q(key_mem[691]), 
	.D(FE_PHN3821_n1555), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_5__50_ (.Q(key_mem[690]), 
	.D(FE_PHN4624_n1556), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_5__49_ (.Q(key_mem[689]), 
	.D(FE_PHN4810_n1557), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_5__44_ (.Q(key_mem[684]), 
	.D(FE_PHN4527_n1562), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_5__43_ (.Q(key_mem[683]), 
	.D(FE_PHN4868_n1563), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_5__41_ (.Q(key_mem[681]), 
	.D(FE_PHN4153_n1565), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_5__39_ (.Q(key_mem[679]), 
	.D(FE_PHN4268_n1567), 
	.CK(clk_48Mhz__L6_N24));
   DFFHQX1 key_mem_reg_5__38_ (.Q(key_mem[678]), 
	.D(FE_PHN4443_n1568), 
	.CK(clk_48Mhz__L6_N3));
   DFFHQX1 key_mem_reg_5__37_ (.Q(key_mem[677]), 
	.D(FE_PHN4642_n1569), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_5__36_ (.Q(key_mem[676]), 
	.D(FE_PHN4625_n1570), 
	.CK(clk_48Mhz__L6_N25));
   DFFHQX1 key_mem_reg_5__35_ (.Q(key_mem[675]), 
	.D(FE_PHN4930_n1571), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 key_mem_reg_5__34_ (.Q(key_mem[674]), 
	.D(FE_PHN4492_n1572), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_5__33_ (.Q(key_mem[673]), 
	.D(FE_PHN4407_n1573), 
	.CK(clk));
   DFFHQX1 key_mem_reg_5__23_ (.Q(key_mem[663]), 
	.D(FE_PHN4613_n1583), 
	.CK(clk_48Mhz__L6_N45));
   DFFHQX1 key_mem_reg_5__22_ (.Q(key_mem[662]), 
	.D(FE_PHN4754_n1584), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_5__21_ (.Q(key_mem[661]), 
	.D(FE_PHN4697_n1585), 
	.CK(clk_48Mhz__L6_N38));
   DFFHQX1 key_mem_reg_5__20_ (.Q(key_mem[660]), 
	.D(FE_PHN4881_n1586), 
	.CK(clk_48Mhz__L6_N42));
   DFFHQX1 key_mem_reg_5__19_ (.Q(key_mem[659]), 
	.D(FE_PHN4803_n1587), 
	.CK(clk_48Mhz__L6_N47));
   DFFHQX1 key_mem_reg_5__18_ (.Q(key_mem[658]), 
	.D(FE_PHN4455_n1588), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_5__17_ (.Q(key_mem[657]), 
	.D(FE_PHN4753_n1589), 
	.CK(clk_48Mhz__L6_N47));
   DFFHQX1 key_mem_reg_5__12_ (.Q(key_mem[652]), 
	.D(FE_PHN3883_n1594), 
	.CK(clk_48Mhz__L6_N18));
   DFFHQX1 key_mem_reg_5__11_ (.Q(key_mem[651]), 
	.D(FE_PHN4446_n1595), 
	.CK(clk_48Mhz__L6_N36));
   DFFHQX1 key_mem_reg_5__9_ (.Q(key_mem[649]), 
	.D(FE_PHN3798_n1597), 
	.CK(clk));
   DFFHQX1 key_mem_reg_5__7_ (.Q(key_mem[647]), 
	.D(FE_PHN4920_n1599), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_5__6_ (.Q(key_mem[646]), 
	.D(FE_PHN916_n1600), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_5__5_ (.Q(key_mem[645]), 
	.D(FE_PHN4748_n1601), 
	.CK(clk_48Mhz__L6_N17));
   DFFHQX1 key_mem_reg_5__4_ (.Q(key_mem[644]), 
	.D(FE_PHN4736_n1602), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_5__3_ (.Q(key_mem[643]), 
	.D(FE_PHN4402_n1603), 
	.CK(clk_48Mhz__L6_N31));
   DFFHQX1 key_mem_reg_5__2_ (.Q(key_mem[642]), 
	.D(FE_PHN3794_n1604), 
	.CK(clk_48Mhz__L6_N14));
   DFFHQX1 key_mem_reg_5__1_ (.Q(key_mem[641]), 
	.D(FE_PHN4781_n1605), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_5__98_ (.Q(key_mem[738]), 
	.D(FE_PHN4905_n1607), 
	.CK(clk_48Mhz__L6_N29));
   DFFHQX1 key_mem_reg_5__97_ (.Q(key_mem[737]), 
	.D(FE_PHN4828_n1608), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_5__87_ (.Q(key_mem[727]), 
	.D(FE_PHN1625_n1618), 
	.CK(clk_48Mhz__L6_N21));
   DFFHQX1 key_mem_reg_5__86_ (.Q(key_mem[726]), 
	.D(FE_PHN4806_n1619), 
	.CK(clk_48Mhz__L6_N33));
   DFFHQX1 key_mem_reg_5__85_ (.Q(key_mem[725]), 
	.D(FE_PHN4200_n1620), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_5__84_ (.Q(key_mem[724]), 
	.D(FE_PHN4927_n1621), 
	.CK(clk_48Mhz__L6_N20));
   DFFHQX1 key_mem_reg_5__83_ (.Q(key_mem[723]), 
	.D(FE_PHN4716_n1622), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_5__82_ (.Q(key_mem[722]), 
	.D(FE_PHN4581_n1623), 
	.CK(clk_48Mhz__L6_N16));
   DFFHQX1 key_mem_reg_5__81_ (.Q(key_mem[721]), 
	.D(FE_PHN4516_n1624), 
	.CK(clk_48Mhz__L6_N7));
   DFFHQX1 key_mem_reg_5__76_ (.Q(key_mem[716]), 
	.D(FE_PHN4735_n1629), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_5__75_ (.Q(key_mem[715]), 
	.D(FE_PHN4833_n1630), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_5__73_ (.Q(key_mem[713]), 
	.D(FE_PHN4825_n1632), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 key_mem_reg_5__71_ (.Q(key_mem[711]), 
	.D(FE_PHN4464_n1634), 
	.CK(clk_48Mhz__L6_N1));
   DFFHQX1 key_mem_reg_5__70_ (.Q(key_mem[710]), 
	.D(FE_PHN4445_n1635), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_5__69_ (.Q(key_mem[709]), 
	.D(FE_PHN4794_n1636), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_5__68_ (.Q(key_mem[708]), 
	.D(FE_PHN4663_n1637), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_5__67_ (.Q(key_mem[707]), 
	.D(FE_PHN4772_n1638), 
	.CK(clk_48Mhz__L6_N32));
   DFFHQX1 key_mem_reg_5__66_ (.Q(key_mem[706]), 
	.D(FE_PHN4574_n1639), 
	.CK(clk_48Mhz__L6_N34));
   DFFHQX1 key_mem_reg_5__65_ (.Q(key_mem[705]), 
	.D(FE_PHN4711_n1640), 
	.CK(clk_48Mhz__L6_N28));
   DFFHQX1 key_mem_reg_5__55_ (.Q(key_mem[695]), 
	.D(FE_PHN4531_n1650), 
	.CK(clk_48Mhz__L6_N13));
   DFFHQX1 key_mem_reg_5__54_ (.Q(key_mem[694]), 
	.D(FE_PHN4776_n1651), 
	.CK(clk_48Mhz__L6_N30));
   DFFHQX1 key_mem_reg_5__53_ (.Q(key_mem[693]), 
	.D(FE_PHN4504_n1652), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_3__119_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1015]), 
	.D(FE_PHN2632_n1277), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_3__118_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1014]), 
	.D(FE_PHN2710_n1278), 
	.CK(clk_48Mhz__L6_N42));
   DFFRHQX1 key_mem_reg_3__117_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1013]), 
	.D(FE_PHN2583_n1279), 
	.CK(clk_48Mhz__L6_N16));
   DFFRHQX1 key_mem_reg_3__116_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1012]), 
	.D(FE_PHN1080_n1280), 
	.CK(clk_48Mhz__L6_N12));
   DFFRHQX1 key_mem_reg_3__115_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1011]), 
	.D(FE_PHN2678_n1281), 
	.CK(clk_48Mhz__L6_N12));
   DFFRHQX1 key_mem_reg_3__114_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1010]), 
	.D(FE_PHN1164_n1282), 
	.CK(clk_48Mhz__L6_N12));
   DFFRHQX1 key_mem_reg_3__113_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1009]), 
	.D(FE_PHN1333_n1283), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_3__108_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1004]), 
	.D(FE_PHN1100_n1288), 
	.CK(clk_48Mhz__L6_N12));
   DFFRHQX1 key_mem_reg_3__107_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1003]), 
	.D(FE_PHN2639_n1289), 
	.CK(clk_48Mhz__L6_N22));
   DFFRHQX1 key_mem_reg_3__105_ (.RN(FE_OFN39_reset_n), 
	.Q(key_mem[1001]), 
	.D(FE_PHN2610_n1291), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 key_mem_reg_3__103_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[999]), 
	.D(FE_PHN2704_n1293), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 key_mem_reg_3__102_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[998]), 
	.D(FE_PHN2775_n1294), 
	.CK(clk_48Mhz__L6_N3));
   DFFRHQX1 key_mem_reg_3__101_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[997]), 
	.D(FE_PHN1088_n1295), 
	.CK(clk_48Mhz__L6_N26));
   DFFRHQX1 key_mem_reg_3__100_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[996]), 
	.D(FE_PHN1092_n1296), 
	.CK(clk_48Mhz__L6_N22));
   DFFRHQX1 key_mem_reg_3__99_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[995]), 
	.D(FE_PHN2539_n1297), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 key_mem_reg_3__98_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[994]), 
	.D(FE_PHN2749_n1298), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 key_mem_reg_3__97_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[993]), 
	.D(FE_PHN1081_n1299), 
	.CK(clk_48Mhz__L6_N34));
   DFFRHQX1 key_mem_reg_3__87_ (.RN(FE_OFN55_reset_n), 
	.Q(key_mem[983]), 
	.D(FE_PHN2615_n1309), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 key_mem_reg_3__86_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[982]), 
	.D(FE_PHN2518_n1310), 
	.CK(clk_48Mhz__L6_N33));
   DFFRHQX1 key_mem_reg_3__85_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[981]), 
	.D(FE_PHN2681_n1311), 
	.CK(clk_48Mhz__L6_N20));
   DFFRHQX1 key_mem_reg_3__84_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[980]), 
	.D(FE_PHN2647_n1312), 
	.CK(clk_48Mhz__L6_N20));
   DFFRHQX1 key_mem_reg_3__83_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[979]), 
	.D(FE_PHN2595_n1313), 
	.CK(clk_48Mhz__L6_N16));
   DFFRHQX1 key_mem_reg_3__82_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[978]), 
	.D(FE_PHN2469_n1314), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 key_mem_reg_3__81_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[977]), 
	.D(FE_PHN2732_n1315), 
	.CK(clk_48Mhz__L6_N7));
   DFFRHQX1 key_mem_reg_3__76_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[972]), 
	.D(FE_PHN995_n1320), 
	.CK(clk_48Mhz__L6_N3));
   DFFRHQX1 key_mem_reg_3__75_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[971]), 
	.D(FE_PHN2593_n1321), 
	.CK(clk_48Mhz__L6_N25));
   DFFRHQX1 key_mem_reg_3__73_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[969]), 
	.D(FE_PHN769_n1323), 
	.CK(clk_48Mhz__L6_N7));
   DFFRHQX1 key_mem_reg_3__71_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[967]), 
	.D(FE_PHN2619_n1325), 
	.CK(clk_48Mhz__L6_N1));
   DFFRHQX1 key_mem_reg_3__70_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[966]), 
	.D(FE_PHN2511_n1326), 
	.CK(clk_48Mhz__L6_N28));
   DFFRHQX1 key_mem_reg_3__69_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[965]), 
	.D(FE_PHN2752_n1327), 
	.CK(clk_48Mhz__L6_N28));
   DFFRHQX1 key_mem_reg_3__68_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[964]), 
	.D(FE_PHN2445_n1328), 
	.CK(clk_48Mhz__L6_N28));
   DFFRHQX1 key_mem_reg_3__67_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[963]), 
	.D(FE_PHN2785_n1329), 
	.CK(clk_48Mhz__L6_N32));
   DFFRHQX1 key_mem_reg_3__66_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[962]), 
	.D(FE_PHN2688_n1330), 
	.CK(clk_48Mhz__L6_N32));
   DFFRHQX1 key_mem_reg_3__65_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[961]), 
	.D(FE_PHN983_n1331), 
	.CK(clk_48Mhz__L6_N28));
   DFFRHQX1 key_mem_reg_3__55_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[951]), 
	.D(FE_PHN2706_n1341), 
	.CK(clk_48Mhz__L6_N13));
   DFFRHQX1 key_mem_reg_3__54_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[950]), 
	.D(FE_PHN796_n1342), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_3__53_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[949]), 
	.D(FE_PHN732_n1343), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_3__52_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[948]), 
	.D(FE_PHN2776_n1344), 
	.CK(clk_48Mhz__L6_N13));
   DFFRHQX1 key_mem_reg_3__51_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[947]), 
	.D(FE_PHN734_n1345), 
	.CK(clk_48Mhz__L6_N17));
   DFFRHQX1 key_mem_reg_3__50_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[946]), 
	.D(FE_PHN2680_n1346), 
	.CK(clk_48Mhz__L6_N13));
   DFFRHQX1 key_mem_reg_3__49_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[945]), 
	.D(FE_PHN2673_n1347), 
	.CK(clk_48Mhz__L6_N24));
   DFFRHQX1 key_mem_reg_3__44_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[940]), 
	.D(FE_PHN2733_n1352), 
	.CK(clk_48Mhz__L6_N31));
   DFFRHQX1 key_mem_reg_3__43_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[939]), 
	.D(FE_PHN2557_n1353), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_3__41_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[937]), 
	.D(FE_PHN2782_n1355), 
	.CK(clk_48Mhz__L6_N28));
   DFFRHQX1 key_mem_reg_3__39_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[935]), 
	.D(FE_PHN2774_n1357), 
	.CK(clk_48Mhz__L6_N24));
   DFFRHQX1 key_mem_reg_3__38_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[934]), 
	.D(FE_PHN2719_n1358), 
	.CK(clk_48Mhz__L6_N3));
   DFFRHQX1 key_mem_reg_3__37_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[933]), 
	.D(FE_PHN2744_n1359), 
	.CK(clk_48Mhz__L6_N28));
   DFFRHQX1 key_mem_reg_3__36_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[932]), 
	.D(FE_PHN733_n1360), 
	.CK(clk_48Mhz__L6_N25));
   DFFRHQX1 key_mem_reg_3__35_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[931]), 
	.D(FE_PHN2763_n1361), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 key_mem_reg_3__34_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[930]), 
	.D(FE_PHN2574_n1362), 
	.CK(clk_48Mhz__L6_N34));
   DFFRHQX1 key_mem_reg_3__33_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[929]), 
	.D(FE_PHN2766_n1363), 
	.CK(clk_48Mhz__L6_N25));
   DFFRHQX1 key_mem_reg_3__23_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[919]), 
	.D(FE_PHN635_n1373), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_3__22_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[918]), 
	.D(FE_PHN2672_n1374), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_3__21_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[917]), 
	.D(FE_PHN2683_n1375), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_3__20_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[916]), 
	.D(FE_PHN998_n1376), 
	.CK(clk_48Mhz__L6_N42));
   DFFRHQX1 key_mem_reg_3__19_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[915]), 
	.D(FE_PHN2708_n1377), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_3__18_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[914]), 
	.D(FE_PHN2714_n1378), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 key_mem_reg_3__17_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[913]), 
	.D(FE_PHN993_n1379), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_3__12_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[908]), 
	.D(FE_PHN2725_n1384), 
	.CK(clk_48Mhz__L6_N18));
   DFFRHQX1 key_mem_reg_3__11_ (.RN(FE_OFN39_reset_n), 
	.Q(key_mem[907]), 
	.D(FE_PHN966_n1385), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 key_mem_reg_3__9_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[905]), 
	.D(FE_PHN2760_n1387), 
	.CK(clk));
   DFFRHQX1 key_mem_reg_3__7_ (.RN(FE_OFN42_reset_n), 
	.Q(key_mem[903]), 
	.D(FE_PHN590_n1389), 
	.CK(clk_48Mhz__L6_N1));
   DFFRHQX1 key_mem_reg_3__6_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[902]), 
	.D(FE_PHN2771_n1390), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 key_mem_reg_3__5_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[901]), 
	.D(FE_PHN988_n1391), 
	.CK(clk_48Mhz__L6_N17));
   DFFRHQX1 key_mem_reg_3__4_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[900]), 
	.D(FE_PHN2715_n1392), 
	.CK(clk_48Mhz__L6_N17));
   DFFRHQX1 key_mem_reg_3__3_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[899]), 
	.D(FE_PHN2781_n1393), 
	.CK(clk_48Mhz__L6_N31));
   DFFRHQX1 key_mem_reg_3__2_ (.RN(FE_OFN55_reset_n), 
	.Q(key_mem[898]), 
	.D(FE_PHN2588_n1394), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 key_mem_reg_3__1_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[897]), 
	.D(FE_PHN948_n1395), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 key_mem_reg_3__121_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1017]), 
	.D(FE_PHN2709_n1275), 
	.CK(clk_48Mhz__L6_N18));
   DFFRHQX1 key_mem_reg_3__89_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[985]), 
	.D(FE_PHN2729_n1307), 
	.CK(clk_48Mhz__L6_N33));
   DFFRHQX1 key_mem_reg_3__57_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[953]), 
	.D(FE_PHN2739_n1339), 
	.CK(clk_48Mhz__L6_N20));
   DFFRHQX1 key_mem_reg_3__25_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[921]), 
	.D(FE_PHN2780_n1371), 
	.CK(clk_48Mhz__L6_N18));
   DFFRHQX1 key_mem_reg_3__123_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1019]), 
	.D(FE_PHN2586_n1273), 
	.CK(clk_48Mhz__L6_N19));
   DFFRHQX1 key_mem_reg_3__91_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[987]), 
	.D(FE_PHN633_n1305), 
	.CK(clk_48Mhz__L6_N16));
   DFFRHQX1 key_mem_reg_3__59_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[955]), 
	.D(FE_PHN2666_n1337), 
	.CK(clk_48Mhz__L6_N17));
   DFFRHQX1 key_mem_reg_3__27_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[923]), 
	.D(FE_PHN2580_n1369), 
	.CK(clk_48Mhz__L6_N18));
   DFFRHQX1 key_mem_reg_3__124_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1020]), 
	.D(FE_PHN2745_n1272), 
	.CK(clk_48Mhz__L6_N12));
   DFFRHQX1 key_mem_reg_3__92_ (.RN(FE_OFN43_reset_n), 
	.Q(key_mem[988]), 
	.D(FE_PHN2643_n1304), 
	.CK(clk_48Mhz__L6_N20));
   DFFRHQX1 key_mem_reg_3__60_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[956]), 
	.D(FE_PHN707_n1336), 
	.CK(clk_48Mhz__L6_N33));
   DFFRHQX1 key_mem_reg_3__28_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[924]), 
	.D(FE_PHN2743_n1368), 
	.CK(clk_48Mhz__L6_N22));
   DFFRHQX1 key_mem_reg_2__119_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1143]), 
	.D(FE_PHN4909_n1149), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_2__118_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1142]), 
	.D(FE_PHN4785_n1150), 
	.CK(clk_48Mhz__L6_N42));
   DFFRHQX1 key_mem_reg_2__117_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1141]), 
	.D(FE_PHN4533_n1151), 
	.CK(clk_48Mhz__L6_N16));
   DFFRHQX1 key_mem_reg_2__116_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1140]), 
	.D(FE_PHN4919_n1152), 
	.CK(clk_48Mhz__L6_N12));
   DFFRHQX1 key_mem_reg_2__115_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1139]), 
	.D(FE_PHN1093_n1153), 
	.CK(clk_48Mhz__L6_N12));
   DFFRHQX1 key_mem_reg_2__114_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1138]), 
	.D(FE_PHN4923_n1154), 
	.CK(clk_48Mhz__L6_N16));
   DFFRHQX1 key_mem_reg_2__113_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1137]), 
	.D(FE_PHN4755_n1155), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 key_mem_reg_2__108_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1132]), 
	.D(FE_PHN4374_n1160), 
	.CK(clk_48Mhz__L6_N16));
   DFFRHQX1 key_mem_reg_2__107_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1131]), 
	.D(FE_PHN428_n1161), 
	.CK(clk_48Mhz__L6_N22));
   DFFRHQX1 key_mem_reg_2__105_ (.RN(FE_OFN39_reset_n), 
	.Q(key_mem[1129]), 
	.D(FE_PHN1323_n1163), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 key_mem_reg_2__103_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1127]), 
	.D(FE_PHN4848_n1165), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 key_mem_reg_2__102_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1126]), 
	.D(FE_PHN1086_n1166), 
	.CK(clk_48Mhz__L6_N1));
   DFFRHQX1 key_mem_reg_2__101_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1125]), 
	.D(FE_PHN1878_n1167), 
	.CK(clk_48Mhz__L6_N26));
   DFFRHQX1 key_mem_reg_2__100_ (.RN(FE_OFN55_reset_n), 
	.Q(key_mem[1124]), 
	.D(FE_PHN1752_n1168), 
	.CK(clk_48Mhz__L6_N26));
   DFFRHQX1 key_mem_reg_2__99_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1123]), 
	.D(FE_PHN4507_n1169), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 key_mem_reg_2__98_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1122]), 
	.D(FE_PHN1098_n1170), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 key_mem_reg_2__97_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1121]), 
	.D(FE_PHN4837_n1171), 
	.CK(clk_48Mhz__L6_N34));
   DFFRHQX1 key_mem_reg_2__87_ (.RN(FE_OFN55_reset_n), 
	.Q(key_mem[1111]), 
	.D(FE_PHN1827_n1181), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 key_mem_reg_2__86_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1110]), 
	.D(FE_PHN999_n1182), 
	.CK(clk_48Mhz__L6_N33));
   DFFRHQX1 key_mem_reg_2__85_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1109]), 
	.D(FE_PHN4686_n1183), 
	.CK(clk_48Mhz__L6_N20));
   DFFRHQX1 key_mem_reg_2__84_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1108]), 
	.D(FE_PHN962_n1184), 
	.CK(clk_48Mhz__L6_N20));
   DFFRHQX1 key_mem_reg_2__83_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1107]), 
	.D(FE_PHN945_n1185), 
	.CK(clk_48Mhz__L6_N16));
   DFFRHQX1 key_mem_reg_2__82_ (.RN(FE_OFN58_reset_n), 
	.Q(key_mem[1106]), 
	.D(FE_PHN4893_n1186), 
	.CK(clk_48Mhz__L6_N16));
   DFFRHQX1 key_mem_reg_2__81_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1105]), 
	.D(FE_PHN4541_n1187), 
	.CK(clk_48Mhz__L6_N7));
   DFFRHQX1 key_mem_reg_2__76_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1100]), 
	.D(FE_PHN4974_n1192), 
	.CK(clk_48Mhz__L6_N3));
   DFFRHQX1 key_mem_reg_2__75_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1099]), 
	.D(FE_PHN4916_n1193), 
	.CK(clk_48Mhz__L6_N25));
   DFFRHQX1 key_mem_reg_2__73_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1097]), 
	.D(FE_PHN4726_n1195), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 key_mem_reg_2__71_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1095]), 
	.D(FE_PHN4500_n1197), 
	.CK(clk_48Mhz__L6_N3));
   DFFRHQX1 key_mem_reg_2__70_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1094]), 
	.D(FE_PHN4891_n1198), 
	.CK(clk_48Mhz__L6_N28));
   DFFRHQX1 key_mem_reg_2__69_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1093]), 
	.D(FE_PHN4820_n1199), 
	.CK(clk_48Mhz__L6_N28));
   DFFRHQX1 key_mem_reg_2__68_ (.RN(FE_OFN40_reset_n), 
	.Q(key_mem[1092]), 
	.D(FE_PHN4750_n1200), 
	.CK(clk_48Mhz__L6_N28));
   DFFRHQX1 key_mem_reg_2__67_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1091]), 
	.D(FE_PHN1016_n1201), 
	.CK(clk_48Mhz__L6_N32));
   DFFRHQX1 key_mem_reg_2__66_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1090]), 
	.D(FE_PHN4758_n1202), 
	.CK(clk_48Mhz__L6_N34));
   DFFRHQX1 key_mem_reg_2__65_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1089]), 
	.D(FE_PHN4850_n1203), 
	.CK(clk_48Mhz__L6_N28));
   DFFRHQX1 key_mem_reg_2__55_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1079]), 
	.D(FE_PHN4766_n1213), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_2__54_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1078]), 
	.D(FE_PHN4902_n1214), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_2__53_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1077]), 
	.D(FE_PHN4733_n1215), 
	.CK(clk_48Mhz__L6_N30));
   DFFRHQX1 key_mem_reg_2__52_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1076]), 
	.D(FE_PHN4757_n1216), 
	.CK(clk_48Mhz__L6_N13));
   DFFRHQX1 key_mem_reg_2__51_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1075]), 
	.D(FE_PHN4372_n1217), 
	.CK(clk_48Mhz__L6_N17));
   DFFRHQX1 key_mem_reg_2__50_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1074]), 
	.D(FE_PHN4401_n1218), 
	.CK(clk_48Mhz__L6_N13));
   DFFRHQX1 key_mem_reg_2__49_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1073]), 
	.D(FE_PHN736_n1219), 
	.CK(clk_48Mhz__L6_N24));
   DFFRHQX1 key_mem_reg_2__44_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1068]), 
	.D(FE_PHN4972_n1224), 
	.CK(clk_48Mhz__L6_N31));
   DFFRHQX1 key_mem_reg_2__43_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1067]), 
	.D(FE_PHN735_n1225), 
	.CK(clk_48Mhz__L6_N31));
   DFFRHQX1 key_mem_reg_2__41_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1065]), 
	.D(FE_PHN1326_n1227), 
	.CK(clk_48Mhz__L6_N24));
   DFFRHQX1 key_mem_reg_2__39_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1063]), 
	.D(FE_PHN4534_n1229), 
	.CK(clk_48Mhz__L6_N24));
   DFFRHQX1 key_mem_reg_2__38_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1062]), 
	.D(FE_PHN2787_n1230), 
	.CK(clk_48Mhz__L6_N3));
   DFFRHQX1 key_mem_reg_2__37_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1061]), 
	.D(FE_PHN4949_n1231), 
	.CK(clk_48Mhz__L6_N25));
   DFFRHQX1 key_mem_reg_2__36_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1060]), 
	.D(FE_PHN4879_n1232), 
	.CK(clk_48Mhz__L6_N25));
   DFFRHQX1 key_mem_reg_2__35_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1059]), 
	.D(FE_PHN4929_n1233), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 key_mem_reg_2__34_ (.RN(FE_OFN36_reset_n), 
	.Q(key_mem[1058]), 
	.D(FE_PHN4485_n1234), 
	.CK(clk_48Mhz__L6_N34));
   DFFRHQX1 key_mem_reg_2__33_ (.RN(FE_OFN37_reset_n), 
	.Q(key_mem[1057]), 
	.D(FE_PHN4672_n1235), 
	.CK(clk));
   DFFRHQX1 key_mem_reg_2__23_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1047]), 
	.D(FE_PHN4555_n1245), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 key_mem_reg_2__22_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1046]), 
	.D(FE_PHN4975_n1246), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_2__21_ (.RN(FE_OFN46_reset_n), 
	.Q(key_mem[1045]), 
	.D(FE_PHN4917_n1247), 
	.CK(clk_48Mhz__L6_N38));
   DFFRHQX1 key_mem_reg_2__20_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1044]), 
	.D(FE_PHN4937_n1248), 
	.CK(clk_48Mhz__L6_N42));
   DFFRHQX1 key_mem_reg_2__19_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1043]), 
	.D(FE_PHN4816_n1249), 
	.CK(clk_48Mhz__L6_N42));
   DFFRHQX1 key_mem_reg_2__18_ (.RN(FE_OFN39_reset_n), 
	.Q(key_mem[1042]), 
	.D(FE_PHN4176_n1250), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 key_mem_reg_2__17_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem[1041]), 
	.D(FE_PHN4842_n1251), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 key_mem_reg_2__12_ (.RN(FE_OFN57_reset_n), 
	.Q(key_mem[1036]), 
	.D(FE_PHN4907_n1256), 
	.CK(clk_48Mhz__L6_N18));
   DFFRHQX1 key_mem_reg_2__11_ (.RN(FE_OFN39_reset_n), 
	.Q(key_mem[1035]), 
	.D(FE_PHN1767_n1257), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 key_mem_reg_2__9_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1033]), 
	.D(FE_PHN588_n1259), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 key_mem_reg_2__7_ (.RN(FE_OFN42_reset_n), 
	.Q(key_mem[1031]), 
	.D(FE_PHN4926_n1261), 
	.CK(clk_48Mhz__L6_N1));
   DFFRHQX1 key_mem_reg_2__6_ (.RN(FE_OFN47_reset_n), 
	.Q(key_mem[1030]), 
	.D(FE_PHN4912_n1262), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 key_mem_reg_2__5_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1029]), 
	.D(FE_PHN4951_n1263), 
	.CK(clk_48Mhz__L6_N17));
   DFFRHQX1 key_mem_reg_2__4_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1028]), 
	.D(FE_PHN4858_n1264), 
	.CK(clk_48Mhz__L6_N17));
   DFFRHQX1 key_mem_reg_2__3_ (.RN(FE_OFN41_reset_n), 
	.Q(key_mem[1027]), 
	.D(FE_PHN996_n1265), 
	.CK(clk_48Mhz__L6_N31));
   DFFRHQX1 key_mem_reg_2__2_ (.RN(FE_OFN55_reset_n), 
	.Q(key_mem[1026]), 
	.D(FE_PHN1774_n1266), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 key_mem_reg_2__1_ (.RN(FE_OFN44_reset_n), 
	.Q(key_mem[1025]), 
	.D(FE_PHN4921_n1267), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 prev_key1_reg_reg_23_ (.Q(FE_PHN1969_keymem_sboxw_23_), 
	.D(FE_PHN5044_n2397), 
	.CK(clk_48Mhz__L6_N37));
   DFFHQX1 prev_key1_reg_reg_15_ (.Q(FE_PHN1972_keymem_sboxw_15_), 
	.D(FE_PHN5039_n2405), 
	.CK(clk_48Mhz__L6_N5));
   DFFHQX1 prev_key1_reg_reg_7_ (.Q(FE_PHN265_keymem_sboxw_7_), 
	.D(FE_PHN5031_n2413), 
	.CK(clk_48Mhz__L6_N2));
   DFFHQX1 prev_key1_reg_reg_31_ (.Q(sboxw[31]), 
	.D(FE_PHN2791_n2389), 
	.CK(clk_48Mhz__L6_N9));
   DFFHQX1 prev_key1_reg_reg_14_ (.Q(FE_PHN1974_keymem_sboxw_14_), 
	.D(FE_PHN5043_n2406), 
	.CK(clk_48Mhz__L6_N5));
   DFFHQX1 prev_key1_reg_reg_30_ (.Q(sboxw[30]), 
	.D(FE_PHN2795_n2390), 
	.CK(clk_48Mhz__L6_N6));
   DFFHQX1 prev_key1_reg_reg_22_ (.Q(sboxw[22]), 
	.D(FE_PHN5041_n2398), 
	.CK(clk_48Mhz__L6_N5));
   DFFHQX1 prev_key1_reg_reg_6_ (.Q(FE_PHN748_keymem_sboxw_6_), 
	.D(FE_PHN5033_n2414), 
	.CK(clk_48Mhz__L6_N5));
   DFFHQX1 prev_key1_reg_reg_26_ (.Q(sboxw[26]), 
	.D(FE_PHN2036_n2394), 
	.CK(clk_48Mhz__L6_N15));
   DFFHQX1 prev_key1_reg_reg_21_ (.Q(sboxw[21]), 
	.D(FE_PHN1463_n2399), 
	.CK(clk_48Mhz__L6_N14));
   DFFHQX1 prev_key1_reg_reg_19_ (.Q(FE_PHN1992_keymem_sboxw_19_), 
	.D(FE_PHN5049_n2401), 
	.CK(clk_48Mhz__L6_N21));
   DFFHQX1 prev_key1_reg_reg_18_ (.Q(sboxw[18]), 
	.D(FE_PHN5037_n2402), 
	.CK(clk_48Mhz__L6_N21));
   DFFHQX1 prev_key1_reg_reg_17_ (.Q(sboxw[17]), 
	.D(FE_PHN5054_n2403), 
	.CK(clk_48Mhz__L6_N11));
   DFFHQX1 prev_key1_reg_reg_16_ (.Q(FE_PHN1997_keymem_sboxw_16_), 
	.D(FE_PHN5051_n2404), 
	.CK(clk_48Mhz__L6_N6));
   DFFHQX1 prev_key1_reg_reg_13_ (.Q(FE_PHN2007_keymem_sboxw_13_), 
	.D(FE_PHN5076_n2407), 
	.CK(clk_48Mhz__L6_N14));
   DFFHQX1 prev_key1_reg_reg_11_ (.Q(FE_PHN2002_keymem_sboxw_11_), 
	.D(FE_PHN5055_n2409), 
	.CK(clk_48Mhz__L6_N14));
   DFFHQX1 prev_key1_reg_reg_10_ (.Q(sboxw[10]), 
	.D(FE_PHN5040_n2410), 
	.CK(clk_48Mhz__L6_N14));
   DFFHQX1 prev_key1_reg_reg_8_ (.Q(sboxw[8]), 
	.D(FE_PHN5056_n2412), 
	.CK(clk_48Mhz__L6_N11));
   DFFHQX1 prev_key1_reg_reg_5_ (.Q(sboxw[5]), 
	.D(FE_PHN5077_n2415), 
	.CK(clk_48Mhz__L6_N23));
   DFFHQX1 prev_key1_reg_reg_3_ (.Q(FE_PHN2000_keymem_sboxw_3_), 
	.D(FE_PHN5052_n2417), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 prev_key1_reg_reg_2_ (.Q(sboxw[2]), 
	.D(FE_PHN1038_n2418), 
	.CK(clk_48Mhz__L6_N35));
   DFFHQX1 prev_key1_reg_reg_1_ (.Q(FE_PHN1957_keymem_sboxw_1_), 
	.D(FE_PHN5035_n2419), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 prev_key1_reg_reg_0_ (.Q(sboxw[0]), 
	.D(FE_PHN5038_n2420), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 prev_key1_reg_reg_25_ (.Q(sboxw[25]), 
	.D(FE_PHN2792_n2395), 
	.CK(clk_48Mhz__L6_N8));
   DFFHQX1 prev_key1_reg_reg_27_ (.Q(sboxw[27]), 
	.D(FE_PHN2038_n2393), 
	.CK(clk_48Mhz__L6_N26));
   DFFHQX1 prev_key1_reg_reg_29_ (.Q(sboxw[29]), 
	.D(FE_PHN2799_n2391), 
	.CK(clk_48Mhz__L6_N14));
   DFFHQX1 prev_key1_reg_reg_24_ (.Q(sboxw[24]), 
	.D(FE_PHN2793_n2396), 
	.CK(clk_48Mhz__L6_N8));
   DFFHQX1 prev_key1_reg_reg_20_ (.Q(sboxw[20]), 
	.D(FE_PHN5063_n2400), 
	.CK(clk_48Mhz__L6_N14));
   DFFHQX1 prev_key1_reg_reg_12_ (.Q(sboxw[12]), 
	.D(FE_PHN5060_n2408), 
	.CK(clk_48Mhz__L6_N14));
   DFFHQX1 prev_key1_reg_reg_9_ (.Q(FE_PHN1991_keymem_sboxw_9_), 
	.D(FE_PHN5050_n2411), 
	.CK(clk_48Mhz__L6_N4));
   DFFHQX1 prev_key1_reg_reg_4_ (.Q(sboxw[4]), 
	.D(FE_PHN5062_n2416), 
	.CK(clk_48Mhz__L6_N23));
   DFFHQX1 prev_key1_reg_reg_28_ (.Q(sboxw[28]), 
	.D(FE_PHN2798_n2392), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 round_ctr_reg_reg_1_ (.RN(FE_OFN39_reset_n), 
	.Q(round_ctr_reg[1]), 
	.D(FE_PHN2855_n2423), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 round_ctr_reg_reg_2_ (.RN(FE_OFN39_reset_n), 
	.Q(round_ctr_reg[2]), 
	.D(FE_PHN2811_n2422), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 round_ctr_reg_reg_3_ (.RN(FE_OFN39_reset_n), 
	.Q(round_ctr_reg[3]), 
	.D(FE_PHN2820_n2421), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 key_mem_ctrl_reg_reg_0_ (.RN(FE_OFN39_reset_n), 
	.Q(key_mem_ctrl_reg[0]), 
	.D(FE_PHN283_n2433), 
	.CK(clk_48Mhz__L6_N36));
   DFFRHQX1 key_mem_ctrl_reg_reg_1_ (.RN(FE_OFN53_reset_n), 
	.Q(key_mem_ctrl_reg[1]), 
	.D(FE_PHN1037_n2432), 
	.CK(clk_48Mhz__L6_N36));
   JKFFRX2 round_ctr_reg_reg_0_ (.RN(FE_OFN39_reset_n), 
	.QN(n6), 
	.Q(round_ctr_reg[0]), 
	.K(n879), 
	.J(FE_PHN155_n3), 
	.CK(clk_48Mhz__L6_N36));
   INVX1 U8 (.Y(n2624), 
	.A(n2699));
   INVX1 U9 (.Y(n2623), 
	.A(n2699));
   INVX1 U10 (.Y(n2622), 
	.A(n2699));
   INVX1 U14 (.Y(n2685), 
	.A(FE_OFN88_n1));
   INVX1 U15 (.Y(n2669), 
	.A(FE_OFN86_n1));
   INVX1 U16 (.Y(n2653), 
	.A(FE_OFN86_n1));
   INVX1 U17 (.Y(n2686), 
	.A(FE_OFN89_n1));
   INVX1 U18 (.Y(n2670), 
	.A(FE_OFN89_n1));
   INVX1 U19 (.Y(n2654), 
	.A(FE_OFN89_n1));
   INVX1 U20 (.Y(n2687), 
	.A(n1));
   INVX1 U21 (.Y(n2671), 
	.A(FE_OFN87_n1));
   INVX1 U22 (.Y(n2655), 
	.A(FE_OFN87_n1));
   INVX1 U23 (.Y(n2688), 
	.A(FE_OFN86_n1));
   INVX1 U24 (.Y(n2672), 
	.A(FE_OFN86_n1));
   INVX1 U25 (.Y(n2656), 
	.A(FE_OFN86_n1));
   INVX1 U26 (.Y(n2699), 
	.A(FE_OFN86_n1));
   INVX1 U27 (.Y(n2698), 
	.A(n1));
   INVX1 U28 (.Y(n2697), 
	.A(FE_OFN88_n1));
   INVX1 U29 (.Y(n2696), 
	.A(FE_OFN86_n1));
   INVX1 U30 (.Y(n2695), 
	.A(n1));
   INVX1 U31 (.Y(n2694), 
	.A(n1));
   INVX1 U32 (.Y(n2693), 
	.A(FE_OFN88_n1));
   INVX1 U33 (.Y(n2692), 
	.A(FE_OFN86_n1));
   INVX1 U34 (.Y(n2691), 
	.A(n1));
   INVX1 U35 (.Y(n2690), 
	.A(n1));
   INVX1 U36 (.Y(n2689), 
	.A(FE_OFN85_n1));
   INVX1 U37 (.Y(n2684), 
	.A(FE_OFN86_n1));
   INVX1 U38 (.Y(n2683), 
	.A(n1));
   INVX1 U39 (.Y(n2682), 
	.A(FE_OFN86_n1));
   INVX1 U40 (.Y(n2681), 
	.A(FE_OFN88_n1));
   INVX1 U41 (.Y(n2680), 
	.A(FE_OFN86_n1));
   INVX1 U42 (.Y(n2679), 
	.A(n1));
   INVX1 U43 (.Y(n2678), 
	.A(FE_OFN89_n1));
   INVX1 U44 (.Y(n2677), 
	.A(FE_OFN88_n1));
   INVX1 U45 (.Y(n2676), 
	.A(FE_OFN86_n1));
   INVX1 U46 (.Y(n2675), 
	.A(FE_OFN87_n1));
   INVX1 U47 (.Y(n2674), 
	.A(FE_OFN89_n1));
   INVX1 U48 (.Y(n2673), 
	.A(n1));
   INVX1 U49 (.Y(n2668), 
	.A(FE_OFN86_n1));
   INVX1 U50 (.Y(n2667), 
	.A(FE_OFN89_n1));
   INVX1 U51 (.Y(n2666), 
	.A(FE_OFN89_n1));
   INVX1 U52 (.Y(n2665), 
	.A(FE_OFN88_n1));
   INVX1 U53 (.Y(n2664), 
	.A(FE_OFN86_n1));
   INVX1 U54 (.Y(n2663), 
	.A(n1));
   INVX1 U55 (.Y(n2662), 
	.A(FE_OFN86_n1));
   INVX1 U56 (.Y(n2661), 
	.A(FE_OFN88_n1));
   INVX1 U57 (.Y(n2660), 
	.A(FE_OFN86_n1));
   INVX1 U58 (.Y(n2659), 
	.A(FE_OFN87_n1));
   INVX1 U59 (.Y(n2658), 
	.A(FE_OFN89_n1));
   INVX1 U60 (.Y(n2657), 
	.A(n1));
   INVX1 U61 (.Y(n2652), 
	.A(FE_OFN86_n1));
   INVX1 U62 (.Y(n2651), 
	.A(FE_OFN89_n1));
   INVX1 U63 (.Y(n2650), 
	.A(FE_OFN89_n1));
   INVX1 U64 (.Y(n2649), 
	.A(FE_OFN88_n1));
   INVX1 U65 (.Y(n2648), 
	.A(FE_OFN86_n1));
   INVX1 U66 (.Y(n2647), 
	.A(n1));
   INVX1 U67 (.Y(n2646), 
	.A(FE_OFN89_n1));
   INVX1 U68 (.Y(n2645), 
	.A(FE_OFN88_n1));
   INVX1 U69 (.Y(n2644), 
	.A(FE_OFN86_n1));
   INVX1 U70 (.Y(n2643), 
	.A(FE_OFN87_n1));
   INVX1 U71 (.Y(n2642), 
	.A(FE_OFN89_n1));
   INVX1 U126 (.Y(n2817), 
	.A(n2));
   INVX2 U131 (.Y(n2818), 
	.A(n2));
   INVX1 U134 (.Y(n2637), 
	.A(FE_OFN88_n1));
   INVX1 U135 (.Y(n2638), 
	.A(FE_OFN89_n1));
   INVX1 U136 (.Y(n2639), 
	.A(FE_OFN87_n1));
   INVX1 U137 (.Y(n2640), 
	.A(FE_OFN86_n1));
   INVX1 U138 (.Y(n2641), 
	.A(n1));
   INVX1 U197 (.Y(n2828), 
	.A(n7));
   INVX1 U201 (.Y(n2824), 
	.A(n7));
   INVX1 U205 (.Y(n2829), 
	.A(n7));
   INVX1 U210 (.Y(n2827), 
	.A(n7));
   INVX1 U212 (.Y(n2784), 
	.A(n5));
   INVX2 U215 (.Y(n2781), 
	.A(n5));
   INVX1 U222 (.Y(n2780), 
	.A(n5));
   INVX1 U225 (.Y(n2769), 
	.A(n4));
   INVX2 U226 (.Y(n2806), 
	.A(n8));
   INVX1 U233 (.Y(n2773), 
	.A(n4));
   INVX1 U235 (.Y(n2770), 
	.A(n4));
   INVX1 U237 (.Y(n2766), 
	.A(n4));
   NOR2XL U306 (.Y(n679), 
	.B(FE_PHN112_round_ctr_reg_1_), 
	.A(n683));
   XOR2X1 U307 (.Y(n731), 
	.B(n765), 
	.A(n692));
   XOR2X1 U308 (.Y(n733), 
	.B(n771), 
	.A(n696));
   XOR2X1 U309 (.Y(n736), 
	.B(n780), 
	.A(n702));
   XOR2X1 U310 (.Y(n738), 
	.B(n786), 
	.A(n706));
   XOR2X1 U311 (.Y(n734), 
	.B(n774), 
	.A(n698));
   XOR2X1 U312 (.Y(n735), 
	.B(n777), 
	.A(n700));
   XOR2X1 U313 (.Y(n737), 
	.B(n783), 
	.A(n704));
   XOR2X1 U314 (.Y(n732), 
	.B(n768), 
	.A(n694));
   OR2X2 U318 (.Y(n1), 
	.B(FE_OFN90_n690), 
	.A(n675));
   INVX4 U320 (.Y(n2823), 
	.A(n7));
   CLKINVX3 U321 (.Y(n2800), 
	.A(n8));
   INVX4 U324 (.Y(n2775), 
	.A(n5));
   OR3XL U329 (.Y(n2), 
	.C(n2878), 
	.B(n2877), 
	.A(n2876));
   NOR2BX4 U330 (.Y(n30), 
	.B(n2876), 
	.AN(n540));
   INVX1 U331 (.Y(n2872), 
	.A(FE_PHN112_round_ctr_reg_1_));
   NAND3BX2 U332 (.Y(n676), 
	.C(n2873), 
	.B(FE_PHN155_n3), 
	.AN(n677));
   OAI221XL U336 (.Y(n2433), 
	.C0(n542), 
	.B1(n2870), 
	.B0(n884), 
	.A1(FE_PHN254_n689), 
	.A0(n675));
   OAI211XL U337 (.Y(n2432), 
	.C0(n675), 
	.B0(n880), 
	.A1(n2871), 
	.A0(n884));
   OAI21XL U338 (.Y(n876), 
	.B0(n2869), 
	.A1(n675), 
	.A0(FE_PHN112_round_ctr_reg_1_));
   NAND2XL U339 (.Y(n879), 
	.B(FE_PHN2814_n880), 
	.A(n675));
   OAI32XL U340 (.Y(n2421), 
	.B1(n2874), 
	.B0(n875), 
	.A2(n677), 
	.A1(n675), 
	.A0(n2873));
   AOI21X1 U341 (.Y(n875), 
	.B0(n876), 
	.A1(n2873), 
	.A0(FE_PHN155_n3));
   NAND2X1 U342 (.Y(n2430), 
	.B(n2875), 
	.A(FE_PHN155_n3));
   OAI2BB2XL U343 (.Y(n1732), 
	.B1(FE_OFN3_n682), 
	.B0(FE_PHN401_n639), 
	.A1N(FE_PHN3410_key_mem_543_), 
	.A0N(FE_OFN3_n682));
   OAI2BB2XL U344 (.Y(n1700), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN423_n607), 
	.A1N(key_mem[575]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U345 (.Y(n1767), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN342_n575), 
	.A1N(key_mem[607]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U346 (.Y(n1653), 
	.B1(FE_OFN3_n682), 
	.B0(FE_PHN622_n543), 
	.A1N(key_mem[639]), 
	.A0N(FE_OFN3_n682));
   OAI2BB2XL U347 (.Y(n1739), 
	.B1(n682), 
	.B0(FE_PHN406_n646), 
	.A1N(key_mem[536]), 
	.A0N(n682));
   OAI2BB2XL U348 (.Y(n1707), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN404_n614), 
	.A1N(key_mem[568]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U349 (.Y(n1774), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN347_n582), 
	.A1N(key_mem[600]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U350 (.Y(n1660), 
	.B1(n682), 
	.B0(FE_PHN568_n550), 
	.A1N(key_mem[632]), 
	.A0N(n682));
   OAI2BB2XL U351 (.Y(n1733), 
	.B1(FE_OFN3_n682), 
	.B0(FE_PHN408_n640), 
	.A1N(key_mem[542]), 
	.A0N(FE_OFN3_n682));
   OAI2BB2XL U352 (.Y(n1701), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN422_n608), 
	.A1N(key_mem[574]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U353 (.Y(n1768), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN344_n576), 
	.A1N(key_mem[606]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U354 (.Y(n1654), 
	.B1(FE_OFN3_n682), 
	.B0(FE_PHN623_n544), 
	.A1N(key_mem[638]), 
	.A0N(FE_OFN3_n682));
   OAI2BB2XL U355 (.Y(n1734), 
	.B1(n682), 
	.B0(FE_PHN400_n641), 
	.A1N(key_mem[541]), 
	.A0N(n682));
   OAI2BB2XL U356 (.Y(n1702), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN393_n609), 
	.A1N(key_mem[573]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U357 (.Y(n1769), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN343_n577), 
	.A1N(key_mem[605]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U358 (.Y(n1655), 
	.B1(n682), 
	.B0(FE_PHN551_n545), 
	.A1N(key_mem[637]), 
	.A0N(n682));
   OAI2BB2XL U359 (.Y(n1735), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN397_n642), 
	.A1N(key_mem[540]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U360 (.Y(n1703), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN392_n610), 
	.A1N(key_mem[572]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U361 (.Y(n1770), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN345_n578), 
	.A1N(key_mem[604]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U362 (.Y(n1656), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN548_n546), 
	.A1N(key_mem[636]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U363 (.Y(n1736), 
	.B1(n682), 
	.B0(FE_PHN399_n643), 
	.A1N(key_mem[539]), 
	.A0N(n682));
   OAI2BB2XL U364 (.Y(n1704), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN386_n611), 
	.A1N(key_mem[571]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U365 (.Y(n1771), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN346_n579), 
	.A1N(key_mem[603]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U366 (.Y(n1657), 
	.B1(n682), 
	.B0(FE_PHN544_n547), 
	.A1N(key_mem[635]), 
	.A0N(n682));
   OAI2BB2XL U367 (.Y(n1737), 
	.B1(n682), 
	.B0(FE_PHN395_n644), 
	.A1N(key_mem[538]), 
	.A0N(n682));
   OAI2BB2XL U368 (.Y(n1705), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN326_n612), 
	.A1N(key_mem[570]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U369 (.Y(n1772), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN547_n580), 
	.A1N(key_mem[602]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U370 (.Y(n1658), 
	.B1(n682), 
	.B0(FE_PHN418_n548), 
	.A1N(key_mem[634]), 
	.A0N(n682));
   OAI2BB2XL U371 (.Y(n1738), 
	.B1(n682), 
	.B0(FE_PHN407_n645), 
	.A1N(key_mem[537]), 
	.A0N(n682));
   OAI2BB2XL U372 (.Y(n1706), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN405_n613), 
	.A1N(key_mem[569]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U373 (.Y(n1773), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN349_n581), 
	.A1N(key_mem[601]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U374 (.Y(n1659), 
	.B1(n682), 
	.B0(FE_PHN567_n549), 
	.A1N(key_mem[633]), 
	.A0N(n682));
   OAI2BB2XL U375 (.Y(n1780), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN543_n588), 
	.A1N(key_mem[594]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U376 (.Y(n1779), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN549_n587), 
	.A1N(key_mem[595]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U377 (.Y(n1778), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN542_n586), 
	.A1N(key_mem[596]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U378 (.Y(n1777), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN539_n585), 
	.A1N(key_mem[597]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U379 (.Y(n1776), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN576_n584), 
	.A1N(key_mem[598]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U380 (.Y(n1775), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN574_n583), 
	.A1N(key_mem[599]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U381 (.Y(n1766), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN609_n574), 
	.A1N(key_mem[608]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U382 (.Y(n1765), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN610_n573), 
	.A1N(key_mem[609]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U383 (.Y(n1764), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN612_n572), 
	.A1N(key_mem[610]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U384 (.Y(n1763), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN553_n670), 
	.A1N(key_mem[512]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U385 (.Y(n1762), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN537_n669), 
	.A1N(key_mem[513]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U386 (.Y(n1761), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN550_n668), 
	.A1N(FE_PHN3437_key_mem_514_), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U387 (.Y(n1760), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN563_n667), 
	.A1N(key_mem[515]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U388 (.Y(n1759), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN562_n666), 
	.A1N(key_mem[516]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U389 (.Y(n1758), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN566_n665), 
	.A1N(key_mem[517]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U390 (.Y(n1757), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN572_n664), 
	.A1N(key_mem[518]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U391 (.Y(n1756), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN324_n663), 
	.A1N(key_mem[519]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U392 (.Y(n1755), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN325_n662), 
	.A1N(key_mem[520]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U393 (.Y(n1754), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN323_n661), 
	.A1N(key_mem[521]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U394 (.Y(n1753), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN541_n660), 
	.A1N(FE_PHN3416_key_mem_522_), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U395 (.Y(n1752), 
	.B1(n682), 
	.B0(FE_PHN554_n659), 
	.A1N(key_mem[523]), 
	.A0N(n682));
   OAI2BB2XL U396 (.Y(n1751), 
	.B1(n682), 
	.B0(FE_PHN560_n658), 
	.A1N(key_mem[524]), 
	.A0N(n682));
   OAI2BB2XL U397 (.Y(n1750), 
	.B1(n682), 
	.B0(FE_PHN552_n657), 
	.A1N(key_mem[525]), 
	.A0N(n682));
   OAI2BB2XL U398 (.Y(n1749), 
	.B1(FE_OFN3_n682), 
	.B0(FE_PHN571_n656), 
	.A1N(key_mem[526]), 
	.A0N(FE_OFN3_n682));
   OAI2BB2XL U399 (.Y(n1748), 
	.B1(FE_OFN3_n682), 
	.B0(FE_PHN327_n655), 
	.A1N(key_mem[527]), 
	.A0N(FE_OFN3_n682));
   OAI2BB2XL U400 (.Y(n1747), 
	.B1(FE_OFN3_n682), 
	.B0(FE_PHN573_n654), 
	.A1N(key_mem[528]), 
	.A0N(FE_OFN3_n682));
   OAI2BB2XL U401 (.Y(n1746), 
	.B1(FE_OFN3_n682), 
	.B0(FE_PHN570_n653), 
	.A1N(key_mem[529]), 
	.A0N(FE_OFN3_n682));
   OAI2BB2XL U402 (.Y(n1745), 
	.B1(n682), 
	.B0(FE_PHN558_n652), 
	.A1N(key_mem[530]), 
	.A0N(n682));
   OAI2BB2XL U403 (.Y(n1744), 
	.B1(FE_OFN3_n682), 
	.B0(FE_PHN569_n651), 
	.A1N(key_mem[531]), 
	.A0N(FE_OFN3_n682));
   OAI2BB2XL U404 (.Y(n1743), 
	.B1(FE_OFN3_n682), 
	.B0(FE_PHN579_n650), 
	.A1N(key_mem[532]), 
	.A0N(FE_OFN3_n682));
   OAI2BB2XL U405 (.Y(n1742), 
	.B1(FE_OFN3_n682), 
	.B0(FE_PHN625_n649), 
	.A1N(key_mem[533]), 
	.A0N(FE_OFN3_n682));
   OAI2BB2XL U406 (.Y(n1741), 
	.B1(FE_OFN3_n682), 
	.B0(FE_PHN564_n648), 
	.A1N(key_mem[534]), 
	.A0N(FE_OFN3_n682));
   OAI2BB2XL U407 (.Y(n1740), 
	.B1(FE_OFN3_n682), 
	.B0(FE_PHN348_n647), 
	.A1N(key_mem[535]), 
	.A0N(FE_OFN3_n682));
   OAI2BB2XL U408 (.Y(n1731), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN383_n638), 
	.A1N(key_mem[544]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U409 (.Y(n1730), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN380_n637), 
	.A1N(key_mem[545]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U410 (.Y(n1729), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN381_n636), 
	.A1N(key_mem[546]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U411 (.Y(n1728), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN379_n635), 
	.A1N(key_mem[547]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U412 (.Y(n1727), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN394_n634), 
	.A1N(key_mem[548]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U413 (.Y(n1726), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN391_n633), 
	.A1N(key_mem[549]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U414 (.Y(n1725), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN396_n632), 
	.A1N(key_mem[550]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U415 (.Y(n1724), 
	.B1(FE_OFN4_n682), 
	.B0(n631), 
	.A1N(key_mem[551]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U416 (.Y(n1723), 
	.B1(FE_OFN4_n682), 
	.B0(n630), 
	.A1N(key_mem[552]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U417 (.Y(n1722), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN705_n629), 
	.A1N(key_mem[553]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U418 (.Y(n1721), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN390_n628), 
	.A1N(key_mem[554]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U419 (.Y(n1720), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN398_n627), 
	.A1N(key_mem[555]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U420 (.Y(n1719), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN388_n626), 
	.A1N(key_mem[556]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U421 (.Y(n1718), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN387_n625), 
	.A1N(key_mem[557]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U422 (.Y(n1717), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN409_n624), 
	.A1N(key_mem[558]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U423 (.Y(n1716), 
	.B1(FE_OFN4_n682), 
	.B0(n623), 
	.A1N(key_mem[559]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U424 (.Y(n1715), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN403_n622), 
	.A1N(key_mem[560]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U425 (.Y(n1714), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN402_n621), 
	.A1N(key_mem[561]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U426 (.Y(n1713), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN384_n620), 
	.A1N(key_mem[562]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U427 (.Y(n1712), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN382_n619), 
	.A1N(key_mem[563]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U428 (.Y(n1711), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN389_n618), 
	.A1N(key_mem[564]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U429 (.Y(n1710), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN385_n617), 
	.A1N(key_mem[565]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U430 (.Y(n1709), 
	.B1(FE_OFN2_n682), 
	.B0(n616), 
	.A1N(key_mem[566]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U431 (.Y(n1708), 
	.B1(FE_OFN2_n682), 
	.B0(n615), 
	.A1N(key_mem[567]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U432 (.Y(n1699), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN540_n606), 
	.A1N(key_mem[576]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U433 (.Y(n1698), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN555_n605), 
	.A1N(key_mem[577]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U434 (.Y(n1697), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN538_n604), 
	.A1N(key_mem[578]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U435 (.Y(n1696), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN546_n603), 
	.A1N(key_mem[579]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U436 (.Y(n1695), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN557_n602), 
	.A1N(key_mem[580]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U437 (.Y(n1694), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN561_n601), 
	.A1N(key_mem[581]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U438 (.Y(n1693), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN578_n600), 
	.A1N(key_mem[582]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U439 (.Y(n1692), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN545_n599), 
	.A1N(key_mem[583]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U440 (.Y(n1691), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN559_n598), 
	.A1N(key_mem[584]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U441 (.Y(n1690), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN416_n597), 
	.A1N(FE_PHN3414_key_mem_585_), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U442 (.Y(n1689), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN565_n596), 
	.A1N(key_mem[586]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U443 (.Y(n1688), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN556_n595), 
	.A1N(key_mem[587]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U444 (.Y(n1687), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN575_n594), 
	.A1N(key_mem[588]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U445 (.Y(n1686), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN577_n593), 
	.A1N(key_mem[589]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U446 (.Y(n1685), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN420_n592), 
	.A1N(key_mem[590]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U447 (.Y(n1684), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN417_n591), 
	.A1N(key_mem[591]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U448 (.Y(n1683), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN421_n590), 
	.A1N(key_mem[592]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U449 (.Y(n1682), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN419_n589), 
	.A1N(key_mem[593]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U450 (.Y(n1681), 
	.B1(FE_OFN4_n682), 
	.B0(FE_PHN606_n571), 
	.A1N(key_mem[611]), 
	.A0N(FE_OFN4_n682));
   OAI2BB2XL U451 (.Y(n1680), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN617_n570), 
	.A1N(key_mem[612]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U452 (.Y(n1679), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN613_n569), 
	.A1N(key_mem[613]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U453 (.Y(n1678), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN605_n568), 
	.A1N(key_mem[614]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U454 (.Y(n1677), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN611_n567), 
	.A1N(key_mem[615]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U455 (.Y(n1676), 
	.B1(FE_OFN5_n682), 
	.B0(FE_PHN607_n566), 
	.A1N(key_mem[616]), 
	.A0N(FE_OFN5_n682));
   OAI2BB2XL U456 (.Y(n1675), 
	.B1(n682), 
	.B0(n565), 
	.A1N(key_mem[617]), 
	.A0N(n682));
   OAI2BB2XL U457 (.Y(n1674), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN608_n564), 
	.A1N(FE_PHN3415_key_mem_618_), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U458 (.Y(n1673), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN615_n563), 
	.A1N(key_mem[619]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U459 (.Y(n1672), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN618_n562), 
	.A1N(key_mem[620]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U460 (.Y(n1671), 
	.B1(n682), 
	.B0(FE_PHN621_n561), 
	.A1N(key_mem[621]), 
	.A0N(n682));
   OAI2BB2XL U461 (.Y(n1670), 
	.B1(FE_OFN3_n682), 
	.B0(n560), 
	.A1N(key_mem[622]), 
	.A0N(FE_OFN3_n682));
   OAI2BB2XL U462 (.Y(n1669), 
	.B1(FE_OFN3_n682), 
	.B0(n559), 
	.A1N(FE_PHN3413_key_mem_623_), 
	.A0N(FE_OFN3_n682));
   OAI2BB2XL U463 (.Y(n1668), 
	.B1(n682), 
	.B0(n558), 
	.A1N(key_mem[624]), 
	.A0N(n682));
   OAI2BB2XL U464 (.Y(n1667), 
	.B1(n682), 
	.B0(n557), 
	.A1N(key_mem[625]), 
	.A0N(n682));
   OAI2BB2XL U465 (.Y(n1666), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN614_n556), 
	.A1N(key_mem[626]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U466 (.Y(n1665), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN619_n555), 
	.A1N(key_mem[627]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U467 (.Y(n1664), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN620_n554), 
	.A1N(key_mem[628]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U468 (.Y(n1663), 
	.B1(FE_OFN2_n682), 
	.B0(FE_PHN616_n553), 
	.A1N(key_mem[629]), 
	.A0N(FE_OFN2_n682));
   OAI2BB2XL U469 (.Y(n1662), 
	.B1(FE_OFN3_n682), 
	.B0(n552), 
	.A1N(key_mem[630]), 
	.A0N(FE_OFN3_n682));
   OAI2BB2XL U470 (.Y(n1661), 
	.B1(FE_OFN3_n682), 
	.B0(FE_PHN624_n551), 
	.A1N(key_mem[631]), 
	.A0N(FE_OFN3_n682));
   OAI2BB2XL U471 (.Y(n1575), 
	.B1(FE_OFN21_n681), 
	.B0(FE_PHN401_n639), 
	.A1N(FE_PHN1706_key_mem_671_), 
	.A0N(FE_OFN21_n681));
   OAI2BB2XL U472 (.Y(n1642), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN423_n607), 
	.A1N(FE_PHN758_key_mem_703_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U473 (.Y(n1610), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN342_n575), 
	.A1N(FE_PHN1596_key_mem_735_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U474 (.Y(n1525), 
	.B1(FE_OFN21_n681), 
	.B0(FE_PHN622_n543), 
	.A1N(FE_PHN762_key_mem_767_), 
	.A0N(FE_OFN21_n681));
   OAI2BB2XL U475 (.Y(n1582), 
	.B1(FE_OFN21_n681), 
	.B0(FE_PHN406_n646), 
	.A1N(FE_PHN1512_key_mem_664_), 
	.A0N(FE_OFN21_n681));
   OAI2BB2XL U476 (.Y(n1649), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN404_n614), 
	.A1N(FE_PHN1771_key_mem_696_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U477 (.Y(n1617), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN347_n582), 
	.A1N(FE_PHN1642_key_mem_728_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U478 (.Y(n1532), 
	.B1(n681), 
	.B0(FE_PHN568_n550), 
	.A1N(FE_PHN772_key_mem_760_), 
	.A0N(n681));
   OAI2BB2XL U479 (.Y(n1576), 
	.B1(FE_OFN21_n681), 
	.B0(FE_PHN408_n640), 
	.A1N(FE_PHN1569_key_mem_670_), 
	.A0N(FE_OFN21_n681));
   OAI2BB2XL U480 (.Y(n1643), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN422_n608), 
	.A1N(FE_PHN1516_key_mem_702_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U481 (.Y(n1611), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN344_n576), 
	.A1N(FE_PHN1680_key_mem_734_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U482 (.Y(n1526), 
	.B1(FE_OFN21_n681), 
	.B0(FE_PHN623_n544), 
	.A1N(FE_PHN756_key_mem_766_), 
	.A0N(FE_OFN21_n681));
   OAI2BB2XL U483 (.Y(n1577), 
	.B1(n681), 
	.B0(FE_PHN400_n641), 
	.A1N(key_mem[669]), 
	.A0N(n681));
   OAI2BB2XL U484 (.Y(n1644), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN393_n609), 
	.A1N(FE_PHN1656_key_mem_701_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U485 (.Y(n1612), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN343_n577), 
	.A1N(FE_PHN1587_key_mem_733_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U486 (.Y(n1527), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN551_n545), 
	.A1N(FE_PHN1602_key_mem_765_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U487 (.Y(n1578), 
	.B1(n681), 
	.B0(FE_PHN397_n642), 
	.A1N(key_mem[668]), 
	.A0N(n681));
   OAI2BB2XL U488 (.Y(n1645), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN392_n610), 
	.A1N(FE_PHN1483_key_mem_700_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U489 (.Y(n1613), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN345_n578), 
	.A1N(FE_PHN1746_key_mem_732_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U490 (.Y(n1528), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN548_n546), 
	.A1N(FE_PHN1765_key_mem_764_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U491 (.Y(n1579), 
	.B1(n681), 
	.B0(FE_PHN399_n643), 
	.A1N(key_mem[667]), 
	.A0N(n681));
   OAI2BB2XL U492 (.Y(n1646), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN386_n611), 
	.A1N(FE_PHN1535_key_mem_699_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U493 (.Y(n1614), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN346_n579), 
	.A1N(FE_PHN1671_key_mem_731_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U494 (.Y(n1529), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN544_n547), 
	.A1N(FE_PHN1552_key_mem_763_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U495 (.Y(n1580), 
	.B1(n681), 
	.B0(FE_PHN395_n644), 
	.A1N(key_mem[666]), 
	.A0N(n681));
   OAI2BB2XL U496 (.Y(n1647), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN326_n612), 
	.A1N(FE_PHN1698_key_mem_698_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U497 (.Y(n1615), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN547_n580), 
	.A1N(FE_PHN1666_key_mem_730_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U498 (.Y(n1530), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN418_n548), 
	.A1N(FE_PHN1531_key_mem_762_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U499 (.Y(n1581), 
	.B1(n681), 
	.B0(FE_PHN407_n645), 
	.A1N(FE_PHN3214_key_mem_665_), 
	.A0N(n681));
   OAI2BB2XL U500 (.Y(n1648), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN405_n613), 
	.A1N(FE_PHN1645_key_mem_697_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U501 (.Y(n1616), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN349_n581), 
	.A1N(FE_PHN1528_key_mem_729_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U502 (.Y(n1531), 
	.B1(n681), 
	.B0(FE_PHN567_n549), 
	.A1N(FE_PHN3196_key_mem_761_), 
	.A0N(n681));
   OAI2BB2XL U503 (.Y(n1652), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN385_n617), 
	.A1N(FE_PHN1731_key_mem_693_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U504 (.Y(n1651), 
	.B1(FE_OFN20_n681), 
	.B0(n616), 
	.A1N(FE_PHN1779_key_mem_694_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U505 (.Y(n1650), 
	.B1(FE_OFN20_n681), 
	.B0(n615), 
	.A1N(FE_PHN939_key_mem_695_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U506 (.Y(n1641), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN540_n606), 
	.A1N(FE_PHN1721_key_mem_704_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U507 (.Y(n1640), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN555_n605), 
	.A1N(FE_PHN1574_key_mem_705_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U508 (.Y(n1639), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN538_n604), 
	.A1N(FE_PHN1561_key_mem_706_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U509 (.Y(n1638), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN546_n603), 
	.A1N(FE_PHN1750_key_mem_707_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U510 (.Y(n1637), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN557_n602), 
	.A1N(FE_PHN1755_key_mem_708_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U511 (.Y(n1636), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN561_n601), 
	.A1N(FE_PHN1794_key_mem_709_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U512 (.Y(n1635), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN578_n600), 
	.A1N(FE_PHN1702_key_mem_710_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U513 (.Y(n1634), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN545_n599), 
	.A1N(FE_PHN1609_key_mem_711_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U514 (.Y(n1633), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN559_n598), 
	.A1N(FE_PHN1524_key_mem_712_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U515 (.Y(n1632), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN416_n597), 
	.A1N(FE_PHN1820_key_mem_713_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U516 (.Y(n1631), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN565_n596), 
	.A1N(FE_PHN1495_key_mem_714_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U517 (.Y(n1630), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN556_n595), 
	.A1N(FE_PHN1678_key_mem_715_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U518 (.Y(n1629), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN575_n594), 
	.A1N(FE_PHN1695_key_mem_716_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U519 (.Y(n1628), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN577_n593), 
	.A1N(FE_PHN1523_key_mem_717_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U520 (.Y(n1627), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN420_n592), 
	.A1N(FE_PHN1521_key_mem_718_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U521 (.Y(n1626), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN417_n591), 
	.A1N(FE_PHN1530_key_mem_719_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U522 (.Y(n1625), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN421_n590), 
	.A1N(FE_PHN1568_key_mem_720_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U523 (.Y(n1624), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN419_n589), 
	.A1N(FE_PHN1718_key_mem_721_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U524 (.Y(n1623), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN543_n588), 
	.A1N(FE_PHN1519_key_mem_722_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U525 (.Y(n1622), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN549_n587), 
	.A1N(FE_PHN1770_key_mem_723_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U526 (.Y(n1621), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN542_n586), 
	.A1N(FE_PHN1831_key_mem_724_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U527 (.Y(n1620), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN539_n585), 
	.A1N(FE_PHN1556_key_mem_725_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U528 (.Y(n1619), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN576_n584), 
	.A1N(FE_PHN1646_key_mem_726_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U529 (.Y(n1618), 
	.B1(n681), 
	.B0(FE_PHN574_n583), 
	.A1N(key_mem[727]), 
	.A0N(n681));
   OAI2BB2XL U530 (.Y(n1609), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN609_n574), 
	.A1N(FE_PHN1520_key_mem_736_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U531 (.Y(n1608), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN610_n573), 
	.A1N(FE_PHN1804_key_mem_737_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U532 (.Y(n1607), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN612_n572), 
	.A1N(FE_PHN1824_key_mem_738_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U533 (.Y(n1606), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN553_n670), 
	.A1N(FE_PHN684_key_mem_640_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U534 (.Y(n1605), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN537_n669), 
	.A1N(FE_PHN683_key_mem_641_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U535 (.Y(n1604), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN550_n668), 
	.A1N(FE_PHN1502_key_mem_642_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U536 (.Y(n1603), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN563_n667), 
	.A1N(FE_PHN1615_key_mem_643_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U537 (.Y(n1602), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN562_n666), 
	.A1N(FE_PHN1809_key_mem_644_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U538 (.Y(n1601), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN566_n665), 
	.A1N(FE_PHN1624_key_mem_645_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U539 (.Y(n1600), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN572_n664), 
	.A1N(key_mem[646]), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U540 (.Y(n1599), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN324_n663), 
	.A1N(FE_PHN1848_key_mem_647_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U541 (.Y(n1598), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN325_n662), 
	.A1N(FE_PHN1722_key_mem_648_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U542 (.Y(n1597), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN323_n661), 
	.A1N(FE_PHN1481_key_mem_649_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U543 (.Y(n1596), 
	.B1(n681), 
	.B0(FE_PHN541_n660), 
	.A1N(FE_PHN2832_key_mem_650_), 
	.A0N(n681));
   OAI2BB2XL U544 (.Y(n1595), 
	.B1(n681), 
	.B0(FE_PHN554_n659), 
	.A1N(key_mem[651]), 
	.A0N(n681));
   OAI2BB2XL U545 (.Y(n1594), 
	.B1(n681), 
	.B0(FE_PHN560_n658), 
	.A1N(FE_PHN914_key_mem_652_), 
	.A0N(n681));
   OAI2BB2XL U546 (.Y(n1593), 
	.B1(n681), 
	.B0(FE_PHN552_n657), 
	.A1N(key_mem[653]), 
	.A0N(n681));
   OAI2BB2XL U547 (.Y(n1592), 
	.B1(FE_OFN21_n681), 
	.B0(FE_PHN571_n656), 
	.A1N(FE_PHN1577_key_mem_654_), 
	.A0N(FE_OFN21_n681));
   OAI2BB2XL U548 (.Y(n1591), 
	.B1(FE_OFN21_n681), 
	.B0(FE_PHN327_n655), 
	.A1N(FE_PHN1588_key_mem_655_), 
	.A0N(FE_OFN21_n681));
   OAI2BB2XL U549 (.Y(n1590), 
	.B1(FE_OFN21_n681), 
	.B0(FE_PHN573_n654), 
	.A1N(FE_PHN1657_key_mem_656_), 
	.A0N(FE_OFN21_n681));
   OAI2BB2XL U550 (.Y(n1589), 
	.B1(FE_OFN21_n681), 
	.B0(FE_PHN570_n653), 
	.A1N(FE_PHN754_key_mem_657_), 
	.A0N(FE_OFN21_n681));
   OAI2BB2XL U551 (.Y(n1588), 
	.B1(FE_OFN21_n681), 
	.B0(FE_PHN558_n652), 
	.A1N(FE_PHN1505_key_mem_658_), 
	.A0N(FE_OFN21_n681));
   OAI2BB2XL U552 (.Y(n1587), 
	.B1(FE_OFN21_n681), 
	.B0(FE_PHN569_n651), 
	.A1N(FE_PHN1744_key_mem_659_), 
	.A0N(FE_OFN21_n681));
   OAI2BB2XL U553 (.Y(n1586), 
	.B1(FE_OFN21_n681), 
	.B0(FE_PHN579_n650), 
	.A1N(FE_PHN1724_key_mem_660_), 
	.A0N(FE_OFN21_n681));
   OAI2BB2XL U554 (.Y(n1585), 
	.B1(FE_OFN21_n681), 
	.B0(FE_PHN625_n649), 
	.A1N(FE_PHN1797_key_mem_661_), 
	.A0N(FE_OFN21_n681));
   OAI2BB2XL U555 (.Y(n1584), 
	.B1(FE_OFN21_n681), 
	.B0(FE_PHN564_n648), 
	.A1N(FE_PHN1687_key_mem_662_), 
	.A0N(FE_OFN21_n681));
   OAI2BB2XL U556 (.Y(n1583), 
	.B1(FE_OFN21_n681), 
	.B0(FE_PHN348_n647), 
	.A1N(FE_PHN1660_key_mem_663_), 
	.A0N(FE_OFN21_n681));
   OAI2BB2XL U557 (.Y(n1574), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN383_n638), 
	.A1N(FE_PHN1581_key_mem_672_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U558 (.Y(n1573), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN380_n637), 
	.A1N(FE_PHN1694_key_mem_673_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U559 (.Y(n1572), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN381_n636), 
	.A1N(FE_PHN1641_key_mem_674_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U560 (.Y(n1571), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN379_n635), 
	.A1N(FE_PHN1749_key_mem_675_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U561 (.Y(n1570), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN394_n634), 
	.A1N(FE_PHN917_key_mem_676_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U562 (.Y(n1569), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN391_n633), 
	.A1N(FE_PHN1661_key_mem_677_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U563 (.Y(n1568), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN396_n632), 
	.A1N(FE_PHN1579_key_mem_678_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U564 (.Y(n1567), 
	.B1(FE_OFN22_n681), 
	.B0(n631), 
	.A1N(FE_PHN1565_key_mem_679_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U565 (.Y(n1566), 
	.B1(FE_OFN22_n681), 
	.B0(n630), 
	.A1N(FE_PHN1696_key_mem_680_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U566 (.Y(n1565), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN705_n629), 
	.A1N(FE_PHN1564_key_mem_681_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U567 (.Y(n1564), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN390_n628), 
	.A1N(FE_PHN1747_key_mem_682_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U568 (.Y(n1563), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN398_n627), 
	.A1N(FE_PHN1575_key_mem_683_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U569 (.Y(n1562), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN388_n626), 
	.A1N(FE_PHN1776_key_mem_684_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U570 (.Y(n1561), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN387_n625), 
	.A1N(FE_PHN1630_key_mem_685_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U571 (.Y(n1560), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN409_n624), 
	.A1N(FE_PHN1593_key_mem_686_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U572 (.Y(n1559), 
	.B1(FE_OFN22_n681), 
	.B0(n623), 
	.A1N(FE_PHN1663_key_mem_687_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U573 (.Y(n1558), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN403_n622), 
	.A1N(FE_PHN1879_key_mem_688_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U574 (.Y(n1557), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN402_n621), 
	.A1N(FE_PHN1763_key_mem_689_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U575 (.Y(n1556), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN384_n620), 
	.A1N(FE_PHN1506_key_mem_690_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U576 (.Y(n1555), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN382_n619), 
	.A1N(FE_PHN1476_key_mem_691_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U577 (.Y(n1554), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN389_n618), 
	.A1N(FE_PHN1638_key_mem_692_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U578 (.Y(n1553), 
	.B1(FE_OFN22_n681), 
	.B0(FE_PHN606_n571), 
	.A1N(FE_PHN1692_key_mem_739_), 
	.A0N(FE_OFN22_n681));
   OAI2BB2XL U579 (.Y(n1552), 
	.B1(n681), 
	.B0(FE_PHN617_n570), 
	.A1N(key_mem[740]), 
	.A0N(n681));
   OAI2BB2XL U580 (.Y(n1551), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN613_n569), 
	.A1N(FE_PHN1606_key_mem_741_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U581 (.Y(n1550), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN605_n568), 
	.A1N(FE_PHN1668_key_mem_742_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U582 (.Y(n1549), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN611_n567), 
	.A1N(FE_PHN580_key_mem_743_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U583 (.Y(n1548), 
	.B1(FE_OFN23_n681), 
	.B0(FE_PHN607_n566), 
	.A1N(FE_PHN1550_key_mem_744_), 
	.A0N(FE_OFN23_n681));
   OAI2BB2XL U584 (.Y(n1547), 
	.B1(n681), 
	.B0(n565), 
	.A1N(key_mem[745]), 
	.A0N(n681));
   OAI2BB2XL U585 (.Y(n1546), 
	.B1(n681), 
	.B0(FE_PHN608_n564), 
	.A1N(FE_PHN3215_key_mem_746_), 
	.A0N(n681));
   OAI2BB2XL U586 (.Y(n1545), 
	.B1(n681), 
	.B0(FE_PHN615_n563), 
	.A1N(key_mem[747]), 
	.A0N(n681));
   OAI2BB2XL U587 (.Y(n1544), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN618_n562), 
	.A1N(FE_PHN1473_key_mem_748_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U588 (.Y(n1543), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN621_n561), 
	.A1N(FE_PHN1500_key_mem_749_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U589 (.Y(n1542), 
	.B1(FE_OFN21_n681), 
	.B0(n560), 
	.A1N(FE_PHN1636_key_mem_750_), 
	.A0N(FE_OFN21_n681));
   OAI2BB2XL U590 (.Y(n1541), 
	.B1(FE_OFN21_n681), 
	.B0(n559), 
	.A1N(FE_PHN1613_key_mem_751_), 
	.A0N(FE_OFN21_n681));
   OAI2BB2XL U591 (.Y(n1540), 
	.B1(FE_OFN21_n681), 
	.B0(n558), 
	.A1N(FE_PHN1590_key_mem_752_), 
	.A0N(FE_OFN21_n681));
   OAI2BB2XL U592 (.Y(n1539), 
	.B1(n681), 
	.B0(n557), 
	.A1N(FE_PHN2824_key_mem_753_), 
	.A0N(n681));
   OAI2BB2XL U593 (.Y(n1538), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN614_n556), 
	.A1N(FE_PHN1536_key_mem_754_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U594 (.Y(n1537), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN619_n555), 
	.A1N(FE_PHN1828_key_mem_755_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U595 (.Y(n1536), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN620_n554), 
	.A1N(FE_PHN1631_key_mem_756_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U596 (.Y(n1535), 
	.B1(FE_OFN20_n681), 
	.B0(FE_PHN616_n553), 
	.A1N(FE_PHN1679_key_mem_757_), 
	.A0N(FE_OFN20_n681));
   OAI2BB2XL U597 (.Y(n1534), 
	.B1(FE_OFN21_n681), 
	.B0(n552), 
	.A1N(FE_PHN1751_key_mem_758_), 
	.A0N(FE_OFN21_n681));
   OAI2BB2XL U598 (.Y(n1533), 
	.B1(FE_OFN21_n681), 
	.B0(FE_PHN624_n551), 
	.A1N(FE_PHN1723_key_mem_759_), 
	.A0N(FE_OFN21_n681));
   INVX1 U599 (.Y(n2870), 
	.A(FE_PHN290_key_mem_ctrl_reg_0_));
   AND2X2 U600 (.Y(n3), 
	.B(FE_PHN120_key_mem_ctrl_reg_1_), 
	.A(n2870));
   INVX1 U601 (.Y(n675), 
	.A(FE_PHN155_n3));
   OAI2BB2XL U602 (.Y(n1889), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN401_n639), 
	.A1N(FE_PHN3184_key_mem_415_), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U603 (.Y(n1857), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN423_n607), 
	.A1N(key_mem[447]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U604 (.Y(n1825), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN342_n575), 
	.A1N(key_mem[479]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U605 (.Y(n1793), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN622_n543), 
	.A1N(FE_PHN3221_key_mem_511_), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U606 (.Y(n1896), 
	.B1(n684), 
	.B0(FE_PHN406_n646), 
	.A1N(key_mem[408]), 
	.A0N(n684));
   OAI2BB2XL U607 (.Y(n1864), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN404_n614), 
	.A1N(key_mem[440]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U608 (.Y(n1832), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN347_n582), 
	.A1N(key_mem[472]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U609 (.Y(n1800), 
	.B1(n684), 
	.B0(FE_PHN568_n550), 
	.A1N(FE_PHN2826_key_mem_504_), 
	.A0N(n684));
   OAI2BB2XL U610 (.Y(n1890), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN408_n640), 
	.A1N(key_mem[414]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U611 (.Y(n1858), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN422_n608), 
	.A1N(key_mem[446]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U612 (.Y(n1826), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN344_n576), 
	.A1N(key_mem[478]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U613 (.Y(n1794), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN623_n544), 
	.A1N(key_mem[510]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U614 (.Y(n1891), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN400_n641), 
	.A1N(key_mem[413]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U615 (.Y(n1859), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN393_n609), 
	.A1N(key_mem[445]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U616 (.Y(n1827), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN343_n577), 
	.A1N(key_mem[477]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U617 (.Y(n1795), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN551_n545), 
	.A1N(key_mem[509]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U618 (.Y(n1892), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN397_n642), 
	.A1N(key_mem[412]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U619 (.Y(n1860), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN392_n610), 
	.A1N(key_mem[444]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U620 (.Y(n1828), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN345_n578), 
	.A1N(key_mem[476]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U621 (.Y(n1796), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN548_n546), 
	.A1N(key_mem[508]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U622 (.Y(n1893), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN399_n643), 
	.A1N(key_mem[411]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U623 (.Y(n1861), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN386_n611), 
	.A1N(key_mem[443]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U624 (.Y(n1829), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN346_n579), 
	.A1N(key_mem[475]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U625 (.Y(n1797), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN544_n547), 
	.A1N(key_mem[507]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U626 (.Y(n1894), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN395_n644), 
	.A1N(key_mem[410]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U627 (.Y(n1862), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN326_n612), 
	.A1N(key_mem[442]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U628 (.Y(n1830), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN547_n580), 
	.A1N(key_mem[474]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U629 (.Y(n1798), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN418_n548), 
	.A1N(key_mem[506]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U630 (.Y(n1895), 
	.B1(n684), 
	.B0(FE_PHN407_n645), 
	.A1N(FE_PHN3425_key_mem_409_), 
	.A0N(n684));
   OAI2BB2XL U631 (.Y(n1863), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN405_n613), 
	.A1N(key_mem[441]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U632 (.Y(n1831), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN349_n581), 
	.A1N(key_mem[473]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U633 (.Y(n1799), 
	.B1(n684), 
	.B0(FE_PHN567_n549), 
	.A1N(key_mem[505]), 
	.A0N(n684));
   OAI2BB2XL U634 (.Y(n1908), 
	.B1(n684), 
	.B0(FE_PHN560_n658), 
	.A1N(key_mem[396]), 
	.A0N(n684));
   OAI2BB2XL U635 (.Y(n1907), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN552_n657), 
	.A1N(key_mem[397]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U636 (.Y(n1906), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN571_n656), 
	.A1N(key_mem[398]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U637 (.Y(n1905), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN327_n655), 
	.A1N(FE_PHN3204_key_mem_399_), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U638 (.Y(n1904), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN573_n654), 
	.A1N(key_mem[400]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U639 (.Y(n1903), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN570_n653), 
	.A1N(key_mem[401]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U640 (.Y(n1902), 
	.B1(n684), 
	.B0(FE_PHN558_n652), 
	.A1N(FE_PHN3195_key_mem_402_), 
	.A0N(n684));
   OAI2BB2XL U641 (.Y(n1901), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN569_n651), 
	.A1N(FE_PHN3218_key_mem_403_), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U642 (.Y(n1900), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN579_n650), 
	.A1N(key_mem[404]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U643 (.Y(n1899), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN625_n649), 
	.A1N(key_mem[405]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U644 (.Y(n1898), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN564_n648), 
	.A1N(key_mem[406]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U645 (.Y(n1897), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN348_n647), 
	.A1N(FE_PHN3209_key_mem_407_), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U646 (.Y(n1888), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN383_n638), 
	.A1N(key_mem[416]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U647 (.Y(n1887), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN380_n637), 
	.A1N(key_mem[417]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U648 (.Y(n1886), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN381_n636), 
	.A1N(key_mem[418]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U649 (.Y(n1885), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN379_n635), 
	.A1N(key_mem[419]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U650 (.Y(n1884), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN394_n634), 
	.A1N(key_mem[420]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U651 (.Y(n1883), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN391_n633), 
	.A1N(key_mem[421]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U652 (.Y(n1882), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN396_n632), 
	.A1N(key_mem[422]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U653 (.Y(n1881), 
	.B1(FE_OFN9_n684), 
	.B0(n631), 
	.A1N(key_mem[423]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U654 (.Y(n1880), 
	.B1(FE_OFN9_n684), 
	.B0(n630), 
	.A1N(key_mem[424]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U655 (.Y(n1879), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN705_n629), 
	.A1N(key_mem[425]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U656 (.Y(n1878), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN390_n628), 
	.A1N(key_mem[426]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U657 (.Y(n1877), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN398_n627), 
	.A1N(key_mem[427]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U658 (.Y(n1876), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN388_n626), 
	.A1N(key_mem[428]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U659 (.Y(n1875), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN387_n625), 
	.A1N(key_mem[429]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U660 (.Y(n1874), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN409_n624), 
	.A1N(key_mem[430]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U661 (.Y(n1873), 
	.B1(FE_OFN9_n684), 
	.B0(n623), 
	.A1N(key_mem[431]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U662 (.Y(n1872), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN403_n622), 
	.A1N(key_mem[432]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U663 (.Y(n1871), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN402_n621), 
	.A1N(key_mem[433]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U664 (.Y(n1870), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN384_n620), 
	.A1N(key_mem[434]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U665 (.Y(n1869), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN382_n619), 
	.A1N(key_mem[435]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U666 (.Y(n1868), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN389_n618), 
	.A1N(key_mem[436]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U667 (.Y(n1867), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN385_n617), 
	.A1N(key_mem[437]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U668 (.Y(n1866), 
	.B1(FE_OFN8_n684), 
	.B0(n616), 
	.A1N(key_mem[438]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U669 (.Y(n1865), 
	.B1(FE_OFN8_n684), 
	.B0(n615), 
	.A1N(key_mem[439]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U670 (.Y(n1856), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN540_n606), 
	.A1N(key_mem[448]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U671 (.Y(n1855), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN555_n605), 
	.A1N(key_mem[449]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U672 (.Y(n1854), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN538_n604), 
	.A1N(key_mem[450]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U673 (.Y(n1853), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN546_n603), 
	.A1N(key_mem[451]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U674 (.Y(n1852), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN557_n602), 
	.A1N(key_mem[452]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U675 (.Y(n1851), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN561_n601), 
	.A1N(key_mem[453]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U676 (.Y(n1850), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN578_n600), 
	.A1N(key_mem[454]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U677 (.Y(n1849), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN545_n599), 
	.A1N(key_mem[455]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U678 (.Y(n1848), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN559_n598), 
	.A1N(key_mem[456]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U679 (.Y(n1847), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN416_n597), 
	.A1N(FE_PHN3197_key_mem_457_), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U680 (.Y(n1846), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN565_n596), 
	.A1N(key_mem[458]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U681 (.Y(n1845), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN556_n595), 
	.A1N(key_mem[459]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U682 (.Y(n1844), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN575_n594), 
	.A1N(key_mem[460]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U683 (.Y(n1843), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN577_n593), 
	.A1N(key_mem[461]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U684 (.Y(n1842), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN420_n592), 
	.A1N(key_mem[462]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U685 (.Y(n1841), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN417_n591), 
	.A1N(key_mem[463]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U686 (.Y(n1840), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN421_n590), 
	.A1N(key_mem[464]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U687 (.Y(n1839), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN419_n589), 
	.A1N(key_mem[465]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U688 (.Y(n1838), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN543_n588), 
	.A1N(key_mem[466]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U689 (.Y(n1837), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN549_n587), 
	.A1N(key_mem[467]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U690 (.Y(n1836), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN542_n586), 
	.A1N(key_mem[468]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U691 (.Y(n1835), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN539_n585), 
	.A1N(key_mem[469]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U692 (.Y(n1834), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN576_n584), 
	.A1N(key_mem[470]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U693 (.Y(n1833), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN574_n583), 
	.A1N(key_mem[471]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U694 (.Y(n1824), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN609_n574), 
	.A1N(key_mem[480]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U695 (.Y(n1823), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN610_n573), 
	.A1N(key_mem[481]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U696 (.Y(n1822), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN612_n572), 
	.A1N(key_mem[482]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U697 (.Y(n1821), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN553_n670), 
	.A1N(key_mem[384]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U698 (.Y(n1820), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN537_n669), 
	.A1N(key_mem[385]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U699 (.Y(n1819), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN550_n668), 
	.A1N(FE_PHN3226_key_mem_386_), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U700 (.Y(n1818), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN563_n667), 
	.A1N(key_mem[387]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U701 (.Y(n1817), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN562_n666), 
	.A1N(key_mem[388]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U702 (.Y(n1816), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN566_n665), 
	.A1N(key_mem[389]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U703 (.Y(n1815), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN572_n664), 
	.A1N(key_mem[390]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U704 (.Y(n1814), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN324_n663), 
	.A1N(key_mem[391]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U705 (.Y(n1813), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN325_n662), 
	.A1N(key_mem[392]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U706 (.Y(n1812), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN323_n661), 
	.A1N(key_mem[393]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U707 (.Y(n1811), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN541_n660), 
	.A1N(FE_PHN3430_key_mem_394_), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U708 (.Y(n1810), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN554_n659), 
	.A1N(key_mem[395]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U709 (.Y(n1809), 
	.B1(FE_OFN6_n684), 
	.B0(n559), 
	.A1N(FE_PHN3213_key_mem_495_), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U710 (.Y(n1808), 
	.B1(n684), 
	.B0(n558), 
	.A1N(key_mem[496]), 
	.A0N(n684));
   OAI2BB2XL U711 (.Y(n1807), 
	.B1(n684), 
	.B0(n557), 
	.A1N(key_mem[497]), 
	.A0N(n684));
   OAI2BB2XL U712 (.Y(n1806), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN614_n556), 
	.A1N(key_mem[498]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U713 (.Y(n1805), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN619_n555), 
	.A1N(key_mem[499]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U714 (.Y(n1804), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN620_n554), 
	.A1N(key_mem[500]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U715 (.Y(n1803), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN616_n553), 
	.A1N(key_mem[501]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U716 (.Y(n1802), 
	.B1(FE_OFN6_n684), 
	.B0(n552), 
	.A1N(key_mem[502]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U717 (.Y(n1801), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN624_n551), 
	.A1N(key_mem[503]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U718 (.Y(n1792), 
	.B1(FE_OFN9_n684), 
	.B0(FE_PHN606_n571), 
	.A1N(key_mem[483]), 
	.A0N(FE_OFN9_n684));
   OAI2BB2XL U719 (.Y(n1791), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN617_n570), 
	.A1N(key_mem[484]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U720 (.Y(n1790), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN613_n569), 
	.A1N(key_mem[485]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U721 (.Y(n1789), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN605_n568), 
	.A1N(key_mem[486]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U722 (.Y(n1788), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN611_n567), 
	.A1N(key_mem[487]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U723 (.Y(n1787), 
	.B1(FE_OFN7_n684), 
	.B0(FE_PHN607_n566), 
	.A1N(key_mem[488]), 
	.A0N(FE_OFN7_n684));
   OAI2BB2XL U724 (.Y(n1786), 
	.B1(n684), 
	.B0(n565), 
	.A1N(key_mem[489]), 
	.A0N(n684));
   OAI2BB2XL U725 (.Y(n1785), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN608_n564), 
	.A1N(FE_PHN3422_key_mem_490_), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U726 (.Y(n1784), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN615_n563), 
	.A1N(key_mem[491]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U727 (.Y(n1783), 
	.B1(FE_OFN8_n684), 
	.B0(FE_PHN618_n562), 
	.A1N(key_mem[492]), 
	.A0N(FE_OFN8_n684));
   OAI2BB2XL U728 (.Y(n1782), 
	.B1(FE_OFN6_n684), 
	.B0(FE_PHN621_n561), 
	.A1N(key_mem[493]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U729 (.Y(n1781), 
	.B1(FE_OFN6_n684), 
	.B0(n560), 
	.A1N(key_mem[494]), 
	.A0N(FE_OFN6_n684));
   OAI2BB2XL U730 (.Y(n2104), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN401_n639), 
	.A1N(FE_PHN3411_key_mem_159_), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U731 (.Y(n1947), 
	.B1(n685), 
	.B0(FE_PHN401_n639), 
	.A1N(FE_PHN764_key_mem_287_), 
	.A0N(n685));
   OAI2BB2XL U732 (.Y(n1517), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN401_n639), 
	.A1N(FE_PHN3210_key_mem_799_), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U733 (.Y(n2072), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN423_n607), 
	.A1N(key_mem[191]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U734 (.Y(n2014), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN423_n607), 
	.A1N(FE_PHN1496_key_mem_319_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U735 (.Y(n1485), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN423_n607), 
	.A1N(key_mem[831]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U736 (.Y(n2139), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN342_n575), 
	.A1N(key_mem[223]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U737 (.Y(n1982), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN342_n575), 
	.A1N(FE_PHN1754_key_mem_351_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U738 (.Y(n1453), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN342_n575), 
	.A1N(FE_PHN3203_key_mem_863_), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U739 (.Y(n2037), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN622_n543), 
	.A1N(FE_PHN3418_key_mem_255_), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U740 (.Y(n1909), 
	.B1(n685), 
	.B0(FE_PHN622_n543), 
	.A1N(FE_PHN1517_key_mem_383_), 
	.A0N(n685));
   OAI2BB2XL U741 (.Y(n1421), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN622_n543), 
	.A1N(FE_PHN3275_key_mem_895_), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U742 (.Y(n2111), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN406_n646), 
	.A1N(key_mem[152]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U743 (.Y(n1954), 
	.B1(n685), 
	.B0(FE_PHN406_n646), 
	.A1N(FE_PHN1634_key_mem_280_), 
	.A0N(n685));
   OAI2BB2XL U744 (.Y(n1524), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN406_n646), 
	.A1N(key_mem[792]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U745 (.Y(n2079), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN404_n614), 
	.A1N(key_mem[184]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U746 (.Y(n2021), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN404_n614), 
	.A1N(FE_PHN1537_key_mem_312_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U747 (.Y(n1492), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN404_n614), 
	.A1N(key_mem[824]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U748 (.Y(n2146), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN347_n582), 
	.A1N(key_mem[216]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U749 (.Y(n1989), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN347_n582), 
	.A1N(FE_PHN1775_key_mem_344_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U750 (.Y(n1460), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN347_n582), 
	.A1N(FE_PHN3207_key_mem_856_), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U751 (.Y(n2044), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN568_n550), 
	.A1N(key_mem[248]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U752 (.Y(n1916), 
	.B1(n685), 
	.B0(FE_PHN568_n550), 
	.A1N(FE_PHN1849_key_mem_376_), 
	.A0N(n685));
   OAI2BB2XL U753 (.Y(n1399), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN568_n550), 
	.A1N(key_mem[888]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U754 (.Y(n2105), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN408_n640), 
	.A1N(key_mem[158]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U755 (.Y(n1948), 
	.B1(n685), 
	.B0(FE_PHN408_n640), 
	.A1N(FE_PHN1477_key_mem_286_), 
	.A0N(n685));
   OAI2BB2XL U756 (.Y(n1518), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN408_n640), 
	.A1N(key_mem[798]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U757 (.Y(n2073), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN422_n608), 
	.A1N(key_mem[190]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U758 (.Y(n2015), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN422_n608), 
	.A1N(FE_PHN1806_key_mem_318_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U759 (.Y(n1486), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN422_n608), 
	.A1N(key_mem[830]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U760 (.Y(n2140), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN344_n576), 
	.A1N(key_mem[222]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U761 (.Y(n1983), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN344_n576), 
	.A1N(FE_PHN1614_key_mem_350_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U762 (.Y(n1454), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN344_n576), 
	.A1N(key_mem[862]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U763 (.Y(n2038), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN623_n544), 
	.A1N(key_mem[254]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U764 (.Y(n1910), 
	.B1(n685), 
	.B0(FE_PHN623_n544), 
	.A1N(FE_PHN1503_key_mem_382_), 
	.A0N(n685));
   OAI2BB2XL U765 (.Y(n1422), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN623_n544), 
	.A1N(key_mem[894]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U766 (.Y(n2106), 
	.B1(n687), 
	.B0(FE_PHN400_n641), 
	.A1N(key_mem[157]), 
	.A0N(n687));
   OAI2BB2XL U767 (.Y(n1949), 
	.B1(n685), 
	.B0(FE_PHN400_n641), 
	.A1N(FE_PHN1802_key_mem_285_), 
	.A0N(n685));
   OAI2BB2XL U768 (.Y(n1519), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN400_n641), 
	.A1N(key_mem[797]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U769 (.Y(n2074), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN393_n609), 
	.A1N(key_mem[189]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U770 (.Y(n2016), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN393_n609), 
	.A1N(FE_PHN1658_key_mem_317_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U771 (.Y(n1487), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN393_n609), 
	.A1N(key_mem[829]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U772 (.Y(n2141), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN343_n577), 
	.A1N(key_mem[221]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U773 (.Y(n1984), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN343_n577), 
	.A1N(FE_PHN1851_key_mem_349_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U774 (.Y(n1455), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN343_n577), 
	.A1N(key_mem[861]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U775 (.Y(n2039), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN551_n545), 
	.A1N(key_mem[253]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U776 (.Y(n1911), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN551_n545), 
	.A1N(FE_PHN1501_key_mem_381_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U777 (.Y(n1423), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN551_n545), 
	.A1N(key_mem[893]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U778 (.Y(n2107), 
	.B1(n687), 
	.B0(FE_PHN397_n642), 
	.A1N(key_mem[156]), 
	.A0N(n687));
   OAI2BB2XL U779 (.Y(n1950), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN397_n642), 
	.A1N(FE_PHN1482_key_mem_284_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U780 (.Y(n1520), 
	.B1(n678), 
	.B0(FE_PHN397_n642), 
	.A1N(key_mem[796]), 
	.A0N(n678));
   OAI2BB2XL U781 (.Y(n2075), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN392_n610), 
	.A1N(key_mem[188]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U782 (.Y(n2017), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN392_n610), 
	.A1N(FE_PHN1710_key_mem_316_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U783 (.Y(n1488), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN392_n610), 
	.A1N(key_mem[828]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U784 (.Y(n2142), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN345_n578), 
	.A1N(key_mem[220]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U785 (.Y(n1985), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN345_n578), 
	.A1N(FE_PHN1725_key_mem_348_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U786 (.Y(n1456), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN345_n578), 
	.A1N(key_mem[860]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U787 (.Y(n2040), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN548_n546), 
	.A1N(key_mem[252]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U788 (.Y(n1912), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN548_n546), 
	.A1N(FE_PHN1670_key_mem_380_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U789 (.Y(n1424), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN548_n546), 
	.A1N(key_mem[892]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U790 (.Y(n2108), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN399_n643), 
	.A1N(key_mem[155]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U791 (.Y(n1951), 
	.B1(n685), 
	.B0(FE_PHN399_n643), 
	.A1N(FE_PHN1518_key_mem_283_), 
	.A0N(n685));
   OAI2BB2XL U792 (.Y(n1521), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN399_n643), 
	.A1N(key_mem[795]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U793 (.Y(n2076), 
	.B1(n687), 
	.B0(FE_PHN386_n611), 
	.A1N(key_mem[187]), 
	.A0N(n687));
   OAI2BB2XL U794 (.Y(n2018), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN386_n611), 
	.A1N(FE_PHN1635_key_mem_315_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U795 (.Y(n1489), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN386_n611), 
	.A1N(key_mem[827]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U796 (.Y(n2143), 
	.B1(n687), 
	.B0(FE_PHN346_n579), 
	.A1N(key_mem[219]), 
	.A0N(n687));
   OAI2BB2XL U797 (.Y(n1986), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN346_n579), 
	.A1N(FE_PHN1572_key_mem_347_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U798 (.Y(n1457), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN346_n579), 
	.A1N(key_mem[859]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U799 (.Y(n2041), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN544_n547), 
	.A1N(key_mem[251]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U800 (.Y(n1913), 
	.B1(n685), 
	.B0(FE_PHN544_n547), 
	.A1N(FE_PHN755_key_mem_379_), 
	.A0N(n685));
   OAI2BB2XL U801 (.Y(n1425), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN544_n547), 
	.A1N(key_mem[891]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U802 (.Y(n2109), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN395_n644), 
	.A1N(key_mem[154]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U803 (.Y(n1952), 
	.B1(n685), 
	.B0(FE_PHN395_n644), 
	.A1N(FE_PHN1554_key_mem_282_), 
	.A0N(n685));
   OAI2BB2XL U804 (.Y(n1522), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN395_n644), 
	.A1N(key_mem[794]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U805 (.Y(n2077), 
	.B1(n687), 
	.B0(FE_PHN326_n612), 
	.A1N(key_mem[186]), 
	.A0N(n687));
   OAI2BB2XL U806 (.Y(n2019), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN326_n612), 
	.A1N(FE_PHN1529_key_mem_314_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U807 (.Y(n1490), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN326_n612), 
	.A1N(key_mem[826]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U808 (.Y(n2144), 
	.B1(n687), 
	.B0(FE_PHN547_n580), 
	.A1N(key_mem[218]), 
	.A0N(n687));
   OAI2BB2XL U809 (.Y(n1987), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN547_n580), 
	.A1N(FE_PHN1690_key_mem_346_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U810 (.Y(n1458), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN547_n580), 
	.A1N(key_mem[858]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U811 (.Y(n2042), 
	.B1(n687), 
	.B0(FE_PHN418_n548), 
	.A1N(key_mem[250]), 
	.A0N(n687));
   OAI2BB2XL U812 (.Y(n1914), 
	.B1(n685), 
	.B0(FE_PHN418_n548), 
	.A1N(FE_PHN1589_key_mem_378_), 
	.A0N(n685));
   OAI2BB2XL U813 (.Y(n1397), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN418_n548), 
	.A1N(key_mem[890]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U814 (.Y(n2110), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN407_n645), 
	.A1N(key_mem[153]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U815 (.Y(n1953), 
	.B1(n685), 
	.B0(FE_PHN407_n645), 
	.A1N(FE_PHN1623_key_mem_281_), 
	.A0N(n685));
   OAI2BB2XL U816 (.Y(n1523), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN407_n645), 
	.A1N(key_mem[793]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U817 (.Y(n2078), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN405_n613), 
	.A1N(key_mem[185]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U818 (.Y(n2020), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN405_n613), 
	.A1N(FE_PHN1584_key_mem_313_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U819 (.Y(n1491), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN405_n613), 
	.A1N(key_mem[825]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U820 (.Y(n2145), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN349_n581), 
	.A1N(key_mem[217]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U821 (.Y(n1988), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN349_n581), 
	.A1N(FE_PHN1739_key_mem_345_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U822 (.Y(n1459), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN349_n581), 
	.A1N(key_mem[857]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U823 (.Y(n2043), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN567_n549), 
	.A1N(key_mem[249]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U824 (.Y(n1915), 
	.B1(n685), 
	.B0(FE_PHN567_n549), 
	.A1N(FE_PHN1515_key_mem_377_), 
	.A0N(n685));
   OAI2BB2XL U825 (.Y(n1398), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN567_n549), 
	.A1N(FE_PHN3270_key_mem_889_), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U826 (.Y(n2164), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN578_n600), 
	.A1N(key_mem[198]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U827 (.Y(n2163), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN545_n599), 
	.A1N(key_mem[199]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U828 (.Y(n2162), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN559_n598), 
	.A1N(key_mem[200]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U829 (.Y(n2161), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN416_n597), 
	.A1N(FE_PHN3424_key_mem_201_), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U830 (.Y(n2160), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN565_n596), 
	.A1N(key_mem[202]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U831 (.Y(n2159), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN556_n595), 
	.A1N(key_mem[203]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U832 (.Y(n2158), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN575_n594), 
	.A1N(key_mem[204]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U833 (.Y(n2157), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN577_n593), 
	.A1N(key_mem[205]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U834 (.Y(n2156), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN420_n592), 
	.A1N(key_mem[206]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U835 (.Y(n2155), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN417_n591), 
	.A1N(key_mem[207]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U836 (.Y(n2154), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN421_n590), 
	.A1N(key_mem[208]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U837 (.Y(n2153), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN419_n589), 
	.A1N(key_mem[209]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U838 (.Y(n2152), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN543_n588), 
	.A1N(key_mem[210]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U839 (.Y(n2151), 
	.B1(n687), 
	.B0(FE_PHN549_n587), 
	.A1N(key_mem[211]), 
	.A0N(n687));
   OAI2BB2XL U840 (.Y(n2150), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN542_n586), 
	.A1N(key_mem[212]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U841 (.Y(n2149), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN539_n585), 
	.A1N(key_mem[213]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U842 (.Y(n2148), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN576_n584), 
	.A1N(key_mem[214]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U843 (.Y(n2147), 
	.B1(n687), 
	.B0(FE_PHN574_n583), 
	.A1N(key_mem[215]), 
	.A0N(n687));
   OAI2BB2XL U844 (.Y(n2138), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN609_n574), 
	.A1N(key_mem[224]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U845 (.Y(n2137), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN610_n573), 
	.A1N(key_mem[225]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U846 (.Y(n2136), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN612_n572), 
	.A1N(key_mem[226]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U847 (.Y(n2135), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN553_n670), 
	.A1N(key_mem[128]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U848 (.Y(n2134), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN537_n669), 
	.A1N(key_mem[129]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U849 (.Y(n2133), 
	.B1(n687), 
	.B0(FE_PHN550_n668), 
	.A1N(FE_PHN3429_key_mem_130_), 
	.A0N(n687));
   OAI2BB2XL U850 (.Y(n2132), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN563_n667), 
	.A1N(key_mem[131]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U851 (.Y(n2131), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN562_n666), 
	.A1N(key_mem[132]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U852 (.Y(n2130), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN566_n665), 
	.A1N(key_mem[133]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U853 (.Y(n2129), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN572_n664), 
	.A1N(key_mem[134]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U854 (.Y(n2128), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN324_n663), 
	.A1N(key_mem[135]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U855 (.Y(n2127), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN325_n662), 
	.A1N(key_mem[136]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U856 (.Y(n2126), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN323_n661), 
	.A1N(key_mem[137]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U857 (.Y(n2125), 
	.B1(n687), 
	.B0(FE_PHN541_n660), 
	.A1N(FE_PHN3428_key_mem_138_), 
	.A0N(n687));
   OAI2BB2XL U858 (.Y(n2124), 
	.B1(n687), 
	.B0(FE_PHN554_n659), 
	.A1N(key_mem[139]), 
	.A0N(n687));
   OAI2BB2XL U859 (.Y(n2123), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN560_n658), 
	.A1N(key_mem[140]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U860 (.Y(n2122), 
	.B1(n687), 
	.B0(FE_PHN552_n657), 
	.A1N(key_mem[141]), 
	.A0N(n687));
   OAI2BB2XL U861 (.Y(n2121), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN571_n656), 
	.A1N(key_mem[142]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U862 (.Y(n2120), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN327_n655), 
	.A1N(FE_PHN3420_key_mem_143_), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U863 (.Y(n2119), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN573_n654), 
	.A1N(key_mem[144]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U864 (.Y(n2118), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN570_n653), 
	.A1N(key_mem[145]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U865 (.Y(n2117), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN558_n652), 
	.A1N(key_mem[146]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U866 (.Y(n2116), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN569_n651), 
	.A1N(key_mem[147]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U867 (.Y(n2115), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN579_n650), 
	.A1N(key_mem[148]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U868 (.Y(n2114), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN625_n649), 
	.A1N(key_mem[149]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U869 (.Y(n2113), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN564_n648), 
	.A1N(key_mem[150]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U870 (.Y(n2112), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN348_n647), 
	.A1N(key_mem[151]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U871 (.Y(n2103), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN383_n638), 
	.A1N(key_mem[160]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U872 (.Y(n2102), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN380_n637), 
	.A1N(key_mem[161]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U873 (.Y(n2101), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN381_n636), 
	.A1N(key_mem[162]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U874 (.Y(n2100), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN379_n635), 
	.A1N(key_mem[163]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U875 (.Y(n2099), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN394_n634), 
	.A1N(key_mem[164]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U876 (.Y(n2098), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN391_n633), 
	.A1N(key_mem[165]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U877 (.Y(n2097), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN396_n632), 
	.A1N(key_mem[166]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U878 (.Y(n2096), 
	.B1(FE_OFN29_n687), 
	.B0(n631), 
	.A1N(key_mem[167]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U879 (.Y(n2095), 
	.B1(FE_OFN29_n687), 
	.B0(n630), 
	.A1N(key_mem[168]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U880 (.Y(n2094), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN705_n629), 
	.A1N(key_mem[169]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U881 (.Y(n2093), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN390_n628), 
	.A1N(key_mem[170]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U882 (.Y(n2092), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN398_n627), 
	.A1N(key_mem[171]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U883 (.Y(n2091), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN388_n626), 
	.A1N(key_mem[172]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U884 (.Y(n2090), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN387_n625), 
	.A1N(key_mem[173]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U885 (.Y(n2089), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN409_n624), 
	.A1N(key_mem[174]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U886 (.Y(n2088), 
	.B1(FE_OFN29_n687), 
	.B0(n623), 
	.A1N(key_mem[175]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U887 (.Y(n2087), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN403_n622), 
	.A1N(key_mem[176]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U888 (.Y(n2086), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN402_n621), 
	.A1N(key_mem[177]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U889 (.Y(n2085), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN384_n620), 
	.A1N(key_mem[178]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U890 (.Y(n2084), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN382_n619), 
	.A1N(key_mem[179]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U891 (.Y(n2083), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN389_n618), 
	.A1N(key_mem[180]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U892 (.Y(n2082), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN385_n617), 
	.A1N(key_mem[181]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U893 (.Y(n2081), 
	.B1(FE_OFN29_n687), 
	.B0(n616), 
	.A1N(key_mem[182]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U894 (.Y(n2080), 
	.B1(FE_OFN29_n687), 
	.B0(n615), 
	.A1N(key_mem[183]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U895 (.Y(n2071), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN540_n606), 
	.A1N(key_mem[192]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U896 (.Y(n2070), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN555_n605), 
	.A1N(key_mem[193]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U897 (.Y(n2069), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN538_n604), 
	.A1N(key_mem[194]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U898 (.Y(n2068), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN546_n603), 
	.A1N(key_mem[195]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U899 (.Y(n2067), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN557_n602), 
	.A1N(key_mem[196]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U900 (.Y(n2066), 
	.B1(FE_OFN29_n687), 
	.B0(FE_PHN561_n601), 
	.A1N(key_mem[197]), 
	.A0N(FE_OFN29_n687));
   OAI2BB2XL U901 (.Y(n2065), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN606_n571), 
	.A1N(key_mem[227]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U902 (.Y(n2064), 
	.B1(n687), 
	.B0(FE_PHN617_n570), 
	.A1N(key_mem[228]), 
	.A0N(n687));
   OAI2BB2XL U903 (.Y(n2063), 
	.B1(n687), 
	.B0(FE_PHN613_n569), 
	.A1N(key_mem[229]), 
	.A0N(n687));
   OAI2BB2XL U904 (.Y(n2062), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN605_n568), 
	.A1N(key_mem[230]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U905 (.Y(n2061), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN611_n567), 
	.A1N(key_mem[231]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U906 (.Y(n2060), 
	.B1(FE_OFN30_n687), 
	.B0(FE_PHN607_n566), 
	.A1N(key_mem[232]), 
	.A0N(FE_OFN30_n687));
   OAI2BB2XL U907 (.Y(n2059), 
	.B1(FE_OFN28_n687), 
	.B0(n565), 
	.A1N(key_mem[233]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U908 (.Y(n2058), 
	.B1(n687), 
	.B0(FE_PHN608_n564), 
	.A1N(FE_PHN3423_key_mem_234_), 
	.A0N(n687));
   OAI2BB2XL U909 (.Y(n2057), 
	.B1(n687), 
	.B0(FE_PHN615_n563), 
	.A1N(key_mem[235]), 
	.A0N(n687));
   OAI2BB2XL U910 (.Y(n2056), 
	.B1(n687), 
	.B0(FE_PHN618_n562), 
	.A1N(key_mem[236]), 
	.A0N(n687));
   OAI2BB2XL U911 (.Y(n2055), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN621_n561), 
	.A1N(key_mem[237]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U912 (.Y(n2054), 
	.B1(FE_OFN28_n687), 
	.B0(n560), 
	.A1N(key_mem[238]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U913 (.Y(n2053), 
	.B1(FE_OFN28_n687), 
	.B0(n559), 
	.A1N(FE_PHN3427_key_mem_239_), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U914 (.Y(n2052), 
	.B1(FE_OFN28_n687), 
	.B0(n558), 
	.A1N(key_mem[240]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U915 (.Y(n2051), 
	.B1(FE_OFN28_n687), 
	.B0(n557), 
	.A1N(key_mem[241]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U916 (.Y(n2050), 
	.B1(n687), 
	.B0(FE_PHN614_n556), 
	.A1N(key_mem[242]), 
	.A0N(n687));
   OAI2BB2XL U917 (.Y(n2049), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN619_n555), 
	.A1N(key_mem[243]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U918 (.Y(n2048), 
	.B1(n687), 
	.B0(FE_PHN620_n554), 
	.A1N(key_mem[244]), 
	.A0N(n687));
   OAI2BB2XL U919 (.Y(n2047), 
	.B1(n687), 
	.B0(FE_PHN616_n553), 
	.A1N(key_mem[245]), 
	.A0N(n687));
   OAI2BB2XL U920 (.Y(n2046), 
	.B1(FE_OFN28_n687), 
	.B0(n552), 
	.A1N(key_mem[246]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U921 (.Y(n2045), 
	.B1(FE_OFN28_n687), 
	.B0(FE_PHN624_n551), 
	.A1N(key_mem[247]), 
	.A0N(FE_OFN28_n687));
   OAI2BB2XL U922 (.Y(n2036), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN705_n629), 
	.A1N(FE_PHN1729_key_mem_297_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U923 (.Y(n2035), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN390_n628), 
	.A1N(FE_PHN1586_key_mem_298_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U924 (.Y(n2034), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN398_n627), 
	.A1N(FE_PHN1545_key_mem_299_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U925 (.Y(n2033), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN388_n626), 
	.A1N(FE_PHN1544_key_mem_300_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U926 (.Y(n2032), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN387_n625), 
	.A1N(FE_PHN1650_key_mem_301_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U927 (.Y(n2031), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN409_n624), 
	.A1N(FE_PHN1785_key_mem_302_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U928 (.Y(n2030), 
	.B1(FE_OFN25_n685), 
	.B0(n623), 
	.A1N(FE_PHN1600_key_mem_303_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U929 (.Y(n2029), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN403_n622), 
	.A1N(FE_PHN1507_key_mem_304_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U930 (.Y(n2028), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN402_n621), 
	.A1N(FE_PHN1557_key_mem_305_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U931 (.Y(n2027), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN384_n620), 
	.A1N(FE_PHN1559_key_mem_306_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U932 (.Y(n2026), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN382_n619), 
	.A1N(FE_PHN1633_key_mem_307_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U933 (.Y(n2025), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN389_n618), 
	.A1N(FE_PHN1691_key_mem_308_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U934 (.Y(n2024), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN385_n617), 
	.A1N(FE_PHN1717_key_mem_309_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U935 (.Y(n2023), 
	.B1(FE_OFN25_n685), 
	.B0(n616), 
	.A1N(FE_PHN1547_key_mem_310_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U936 (.Y(n2022), 
	.B1(FE_OFN26_n685), 
	.B0(n615), 
	.A1N(FE_PHN1795_key_mem_311_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U937 (.Y(n2013), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN540_n606), 
	.A1N(FE_PHN1555_key_mem_320_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U938 (.Y(n2012), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN555_n605), 
	.A1N(FE_PHN1621_key_mem_321_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U939 (.Y(n2011), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN538_n604), 
	.A1N(FE_PHN1667_key_mem_322_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U940 (.Y(n2010), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN546_n603), 
	.A1N(FE_PHN1683_key_mem_323_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U941 (.Y(n2009), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN557_n602), 
	.A1N(FE_PHN1716_key_mem_324_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U942 (.Y(n2008), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN561_n601), 
	.A1N(FE_PHN1689_key_mem_325_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U943 (.Y(n2007), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN578_n600), 
	.A1N(FE_PHN1479_key_mem_326_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U944 (.Y(n2006), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN545_n599), 
	.A1N(FE_PHN1543_key_mem_327_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U945 (.Y(n2005), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN559_n598), 
	.A1N(FE_PHN1742_key_mem_328_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U946 (.Y(n2004), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN416_n597), 
	.A1N(FE_PHN1627_key_mem_329_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U947 (.Y(n2003), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN565_n596), 
	.A1N(FE_PHN1603_key_mem_330_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U948 (.Y(n2002), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN556_n595), 
	.A1N(FE_PHN1475_key_mem_331_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U949 (.Y(n2001), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN575_n594), 
	.A1N(FE_PHN1514_key_mem_332_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U950 (.Y(n2000), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN577_n593), 
	.A1N(FE_PHN1472_key_mem_333_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U951 (.Y(n1999), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN420_n592), 
	.A1N(FE_PHN1826_key_mem_334_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U952 (.Y(n1998), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN417_n591), 
	.A1N(FE_PHN1494_key_mem_335_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U953 (.Y(n1997), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN421_n590), 
	.A1N(FE_PHN1493_key_mem_336_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U954 (.Y(n1996), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN419_n589), 
	.A1N(FE_PHN1533_key_mem_337_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U955 (.Y(n1995), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN543_n588), 
	.A1N(FE_PHN1637_key_mem_338_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U956 (.Y(n1994), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN549_n587), 
	.A1N(FE_PHN1464_key_mem_339_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U957 (.Y(n1993), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN542_n586), 
	.A1N(FE_PHN1620_key_mem_340_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U958 (.Y(n1992), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN539_n585), 
	.A1N(FE_PHN1714_key_mem_341_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U959 (.Y(n1991), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN576_n584), 
	.A1N(FE_PHN1653_key_mem_342_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U960 (.Y(n1990), 
	.B1(FE_OFN24_n685), 
	.B0(FE_PHN574_n583), 
	.A1N(FE_PHN1707_key_mem_343_), 
	.A0N(FE_OFN24_n685));
   OAI2BB2XL U961 (.Y(n1981), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN609_n574), 
	.A1N(FE_PHN1844_key_mem_352_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U962 (.Y(n1980), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN610_n573), 
	.A1N(FE_PHN1793_key_mem_353_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U963 (.Y(n1979), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN612_n572), 
	.A1N(FE_PHN1659_key_mem_354_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U964 (.Y(n1978), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN553_n670), 
	.A1N(FE_PHN1711_key_mem_256_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U965 (.Y(n1977), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN537_n669), 
	.A1N(FE_PHN1553_key_mem_257_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U966 (.Y(n1976), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN550_n668), 
	.A1N(FE_PHN1703_key_mem_258_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U967 (.Y(n1975), 
	.B1(FE_OFN25_n685), 
	.B0(FE_PHN563_n667), 
	.A1N(FE_PHN1546_key_mem_259_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U968 (.Y(n1974), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN562_n666), 
	.A1N(FE_PHN1738_key_mem_260_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U969 (.Y(n1973), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN566_n665), 
	.A1N(FE_PHN1652_key_mem_261_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U970 (.Y(n1972), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN572_n664), 
	.A1N(FE_PHN1699_key_mem_262_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U971 (.Y(n1971), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN324_n663), 
	.A1N(FE_PHN1682_key_mem_263_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U972 (.Y(n1970), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN325_n662), 
	.A1N(FE_PHN1632_key_mem_264_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U973 (.Y(n1969), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN323_n661), 
	.A1N(FE_PHN1688_key_mem_265_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U974 (.Y(n1968), 
	.B1(FE_OFN24_n685), 
	.B0(FE_PHN541_n660), 
	.A1N(FE_PHN1697_key_mem_266_), 
	.A0N(FE_OFN24_n685));
   OAI2BB2XL U975 (.Y(n1967), 
	.B1(n685), 
	.B0(FE_PHN554_n659), 
	.A1N(key_mem[267]), 
	.A0N(n685));
   OAI2BB2XL U976 (.Y(n1966), 
	.B1(n685), 
	.B0(FE_PHN560_n658), 
	.A1N(FE_PHN1571_key_mem_268_), 
	.A0N(n685));
   OAI2BB2XL U977 (.Y(n1965), 
	.B1(n685), 
	.B0(FE_PHN552_n657), 
	.A1N(FE_PHN1727_key_mem_269_), 
	.A0N(n685));
   OAI2BB2XL U978 (.Y(n1964), 
	.B1(n685), 
	.B0(FE_PHN571_n656), 
	.A1N(FE_PHN1626_key_mem_270_), 
	.A0N(n685));
   OAI2BB2XL U979 (.Y(n1963), 
	.B1(n685), 
	.B0(FE_PHN327_n655), 
	.A1N(FE_PHN1504_key_mem_271_), 
	.A0N(n685));
   OAI2BB2XL U980 (.Y(n1962), 
	.B1(n685), 
	.B0(FE_PHN573_n654), 
	.A1N(FE_PHN1672_key_mem_272_), 
	.A0N(n685));
   OAI2BB2XL U981 (.Y(n1961), 
	.B1(n685), 
	.B0(FE_PHN570_n653), 
	.A1N(FE_PHN1542_key_mem_273_), 
	.A0N(n685));
   OAI2BB2XL U982 (.Y(n1960), 
	.B1(n685), 
	.B0(FE_PHN558_n652), 
	.A1N(FE_PHN1639_key_mem_274_), 
	.A0N(n685));
   OAI2BB2XL U983 (.Y(n1959), 
	.B1(n685), 
	.B0(FE_PHN569_n651), 
	.A1N(FE_PHN763_key_mem_275_), 
	.A0N(n685));
   OAI2BB2XL U984 (.Y(n1958), 
	.B1(n685), 
	.B0(FE_PHN579_n650), 
	.A1N(FE_PHN1522_key_mem_276_), 
	.A0N(n685));
   OAI2BB2XL U985 (.Y(n1957), 
	.B1(n685), 
	.B0(FE_PHN625_n649), 
	.A1N(FE_PHN1484_key_mem_277_), 
	.A0N(n685));
   OAI2BB2XL U986 (.Y(n1956), 
	.B1(n685), 
	.B0(FE_PHN564_n648), 
	.A1N(FE_PHN1622_key_mem_278_), 
	.A0N(n685));
   OAI2BB2XL U987 (.Y(n1955), 
	.B1(n685), 
	.B0(FE_PHN348_n647), 
	.A1N(FE_PHN1715_key_mem_279_), 
	.A0N(n685));
   OAI2BB2XL U988 (.Y(n1946), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN383_n638), 
	.A1N(FE_PHN1684_key_mem_288_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U989 (.Y(n1945), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN380_n637), 
	.A1N(FE_PHN1492_key_mem_289_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U990 (.Y(n1944), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN381_n636), 
	.A1N(FE_PHN1573_key_mem_290_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U991 (.Y(n1943), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN379_n635), 
	.A1N(FE_PHN1735_key_mem_291_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U992 (.Y(n1942), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN394_n634), 
	.A1N(FE_PHN1525_key_mem_292_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U993 (.Y(n1941), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN391_n633), 
	.A1N(FE_PHN1616_key_mem_293_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U994 (.Y(n1940), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN396_n632), 
	.A1N(FE_PHN1601_key_mem_294_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U995 (.Y(n1939), 
	.B1(FE_OFN25_n685), 
	.B0(n631), 
	.A1N(FE_PHN1511_key_mem_295_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U996 (.Y(n1938), 
	.B1(FE_OFN25_n685), 
	.B0(n630), 
	.A1N(FE_PHN1562_key_mem_296_), 
	.A0N(FE_OFN25_n685));
   OAI2BB2XL U997 (.Y(n1937), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN606_n571), 
	.A1N(FE_PHN1619_key_mem_355_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U998 (.Y(n1936), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN617_n570), 
	.A1N(FE_PHN1549_key_mem_356_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U999 (.Y(n1935), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN613_n569), 
	.A1N(FE_PHN1583_key_mem_357_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U1000 (.Y(n1934), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN605_n568), 
	.A1N(FE_PHN1655_key_mem_358_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U1001 (.Y(n1933), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN611_n567), 
	.A1N(FE_PHN1757_key_mem_359_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U1002 (.Y(n1932), 
	.B1(FE_OFN27_n685), 
	.B0(FE_PHN607_n566), 
	.A1N(FE_PHN1807_key_mem_360_), 
	.A0N(FE_OFN27_n685));
   OAI2BB2XL U1003 (.Y(n1931), 
	.B1(n685), 
	.B0(n565), 
	.A1N(FE_PHN1595_key_mem_361_), 
	.A0N(n685));
   OAI2BB2XL U1004 (.Y(n1930), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN608_n564), 
	.A1N(FE_PHN1594_key_mem_362_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U1005 (.Y(n1929), 
	.B1(FE_OFN24_n685), 
	.B0(FE_PHN615_n563), 
	.A1N(FE_PHN1677_key_mem_363_), 
	.A0N(FE_OFN24_n685));
   OAI2BB2XL U1006 (.Y(n1928), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN618_n562), 
	.A1N(FE_PHN1607_key_mem_364_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U1007 (.Y(n1927), 
	.B1(n685), 
	.B0(FE_PHN621_n561), 
	.A1N(FE_PHN1618_key_mem_365_), 
	.A0N(n685));
   OAI2BB2XL U1008 (.Y(n1926), 
	.B1(n685), 
	.B0(n560), 
	.A1N(FE_PHN1538_key_mem_366_), 
	.A0N(n685));
   OAI2BB2XL U1009 (.Y(n1925), 
	.B1(n685), 
	.B0(n559), 
	.A1N(FE_PHN424_key_mem_367_), 
	.A0N(n685));
   OAI2BB2XL U1010 (.Y(n1924), 
	.B1(n685), 
	.B0(n558), 
	.A1N(FE_PHN1563_key_mem_368_), 
	.A0N(n685));
   OAI2BB2XL U1011 (.Y(n1923), 
	.B1(n685), 
	.B0(n557), 
	.A1N(FE_PHN1605_key_mem_369_), 
	.A0N(n685));
   OAI2BB2XL U1012 (.Y(n1922), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN614_n556), 
	.A1N(FE_PHN1644_key_mem_370_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U1013 (.Y(n1921), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN619_n555), 
	.A1N(FE_PHN915_key_mem_371_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U1014 (.Y(n1920), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN620_n554), 
	.A1N(FE_PHN1580_key_mem_372_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U1015 (.Y(n1919), 
	.B1(FE_OFN26_n685), 
	.B0(FE_PHN616_n553), 
	.A1N(FE_PHN1498_key_mem_373_), 
	.A0N(FE_OFN26_n685));
   OAI2BB2XL U1016 (.Y(n1918), 
	.B1(n685), 
	.B0(n552), 
	.A1N(FE_PHN1726_key_mem_374_), 
	.A0N(n685));
   OAI2BB2XL U1017 (.Y(n1917), 
	.B1(n685), 
	.B0(FE_PHN624_n551), 
	.A1N(FE_PHN1598_key_mem_375_), 
	.A0N(n685));
   OAI2BB2XL U1018 (.Y(n1516), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN383_n638), 
	.A1N(key_mem[800]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1019 (.Y(n1515), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN380_n637), 
	.A1N(key_mem[801]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1020 (.Y(n1514), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN381_n636), 
	.A1N(key_mem[802]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1021 (.Y(n1513), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN379_n635), 
	.A1N(key_mem[803]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1022 (.Y(n1512), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN394_n634), 
	.A1N(key_mem[804]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1023 (.Y(n1511), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN391_n633), 
	.A1N(key_mem[805]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1024 (.Y(n1510), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN396_n632), 
	.A1N(FE_PHN1532_key_mem_806_), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1025 (.Y(n1509), 
	.B1(FE_OFN18_n678), 
	.B0(n631), 
	.A1N(key_mem[807]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1026 (.Y(n1508), 
	.B1(FE_OFN18_n678), 
	.B0(n630), 
	.A1N(key_mem[808]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1027 (.Y(n1507), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN705_n629), 
	.A1N(key_mem[809]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1028 (.Y(n1506), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN390_n628), 
	.A1N(key_mem[810]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U1029 (.Y(n1505), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN398_n627), 
	.A1N(FE_PHN1560_key_mem_811_), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U1030 (.Y(n1504), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN388_n626), 
	.A1N(key_mem[812]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1031 (.Y(n1503), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN387_n625), 
	.A1N(key_mem[813]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1032 (.Y(n1502), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN409_n624), 
	.A1N(key_mem[814]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1033 (.Y(n1501), 
	.B1(FE_OFN18_n678), 
	.B0(n623), 
	.A1N(key_mem[815]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1034 (.Y(n1500), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN403_n622), 
	.A1N(key_mem[816]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1035 (.Y(n1499), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN402_n621), 
	.A1N(key_mem[817]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1036 (.Y(n1498), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN384_n620), 
	.A1N(key_mem[818]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U1037 (.Y(n1497), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN382_n619), 
	.A1N(key_mem[819]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U1038 (.Y(n1496), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN389_n618), 
	.A1N(key_mem[820]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U1039 (.Y(n1495), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN385_n617), 
	.A1N(key_mem[821]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U1040 (.Y(n1494), 
	.B1(FE_OFN17_n678), 
	.B0(n616), 
	.A1N(key_mem[822]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U1041 (.Y(n1493), 
	.B1(FE_OFN17_n678), 
	.B0(n615), 
	.A1N(key_mem[823]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U1042 (.Y(n1484), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN540_n606), 
	.A1N(key_mem[832]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1043 (.Y(n1483), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN555_n605), 
	.A1N(key_mem[833]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1044 (.Y(n1482), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN538_n604), 
	.A1N(key_mem[834]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1045 (.Y(n1481), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN546_n603), 
	.A1N(FE_PHN1469_key_mem_835_), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1046 (.Y(n1480), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN557_n602), 
	.A1N(key_mem[836]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1047 (.Y(n1479), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN561_n601), 
	.A1N(key_mem[837]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1048 (.Y(n1478), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN578_n600), 
	.A1N(key_mem[838]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1049 (.Y(n1477), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN545_n599), 
	.A1N(key_mem[839]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1050 (.Y(n1476), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN559_n598), 
	.A1N(FE_PHN1491_key_mem_840_), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1051 (.Y(n1475), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN416_n597), 
	.A1N(FE_PHN3186_key_mem_841_), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1052 (.Y(n1474), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN565_n596), 
	.A1N(key_mem[842]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1053 (.Y(n1473), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN556_n595), 
	.A1N(key_mem[843]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1054 (.Y(n1472), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN575_n594), 
	.A1N(key_mem[844]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1055 (.Y(n1471), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN577_n593), 
	.A1N(key_mem[845]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1056 (.Y(n1470), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN420_n592), 
	.A1N(FE_PHN2789_key_mem_846_), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1057 (.Y(n1469), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN417_n591), 
	.A1N(key_mem[847]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1058 (.Y(n1468), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN421_n590), 
	.A1N(key_mem[848]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1059 (.Y(n1467), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN419_n589), 
	.A1N(key_mem[849]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1060 (.Y(n1466), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN543_n588), 
	.A1N(key_mem[850]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U1061 (.Y(n1465), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN549_n587), 
	.A1N(key_mem[851]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U1062 (.Y(n1464), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN542_n586), 
	.A1N(key_mem[852]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U1063 (.Y(n1463), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN539_n585), 
	.A1N(key_mem[853]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U1064 (.Y(n1462), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN576_n584), 
	.A1N(key_mem[854]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U1065 (.Y(n1461), 
	.B1(n678), 
	.B0(FE_PHN574_n583), 
	.A1N(key_mem[855]), 
	.A0N(n678));
   OAI2BB2XL U1066 (.Y(n1452), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN609_n574), 
	.A1N(key_mem[864]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1067 (.Y(n1451), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN610_n573), 
	.A1N(key_mem[865]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1068 (.Y(n1450), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN612_n572), 
	.A1N(key_mem[866]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U1069 (.Y(n1449), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN553_n670), 
	.A1N(key_mem[768]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1070 (.Y(n1448), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN537_n669), 
	.A1N(key_mem[769]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1071 (.Y(n1447), 
	.B1(n678), 
	.B0(FE_PHN550_n668), 
	.A1N(FE_PHN3412_key_mem_770_), 
	.A0N(n678));
   OAI2BB2XL U1072 (.Y(n1446), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN563_n667), 
	.A1N(key_mem[771]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1073 (.Y(n1445), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN562_n666), 
	.A1N(key_mem[772]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U1074 (.Y(n1444), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN566_n665), 
	.A1N(key_mem[773]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U1075 (.Y(n1443), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN572_n664), 
	.A1N(key_mem[774]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1076 (.Y(n1442), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN324_n663), 
	.A1N(key_mem[775]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1077 (.Y(n1441), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN325_n662), 
	.A1N(key_mem[776]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1078 (.Y(n1440), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN323_n661), 
	.A1N(FE_PHN3417_key_mem_777_), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1079 (.Y(n1439), 
	.B1(n678), 
	.B0(FE_PHN541_n660), 
	.A1N(key_mem[778]), 
	.A0N(n678));
   OAI2BB2XL U1080 (.Y(n1438), 
	.B1(n678), 
	.B0(FE_PHN554_n659), 
	.A1N(key_mem[779]), 
	.A0N(n678));
   OAI2BB2XL U1081 (.Y(n1437), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN560_n658), 
	.A1N(key_mem[780]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U1082 (.Y(n1436), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN552_n657), 
	.A1N(key_mem[781]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1083 (.Y(n1435), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN571_n656), 
	.A1N(key_mem[782]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U1084 (.Y(n1434), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN327_n655), 
	.A1N(FE_PHN3234_key_mem_783_), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U1085 (.Y(n1433), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN573_n654), 
	.A1N(key_mem[784]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U1086 (.Y(n1432), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN570_n653), 
	.A1N(key_mem[785]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U1087 (.Y(n1431), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN558_n652), 
	.A1N(key_mem[786]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U1088 (.Y(n1430), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN569_n651), 
	.A1N(key_mem[787]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U1089 (.Y(n1429), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN579_n650), 
	.A1N(key_mem[788]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U1090 (.Y(n1428), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN625_n649), 
	.A1N(key_mem[789]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U1091 (.Y(n1427), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN564_n648), 
	.A1N(key_mem[790]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U1092 (.Y(n1426), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN348_n647), 
	.A1N(FE_PHN3198_key_mem_791_), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U1093 (.Y(n1420), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN606_n571), 
	.A1N(key_mem[867]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1094 (.Y(n1419), 
	.B1(n678), 
	.B0(FE_PHN617_n570), 
	.A1N(key_mem[868]), 
	.A0N(n678));
   OAI2BB2XL U1095 (.Y(n1418), 
	.B1(n678), 
	.B0(FE_PHN613_n569), 
	.A1N(key_mem[869]), 
	.A0N(n678));
   OAI2BB2XL U1096 (.Y(n1417), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN605_n568), 
	.A1N(key_mem[870]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1097 (.Y(n1416), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN611_n567), 
	.A1N(key_mem[871]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1098 (.Y(n1415), 
	.B1(FE_OFN18_n678), 
	.B0(FE_PHN607_n566), 
	.A1N(key_mem[872]), 
	.A0N(FE_OFN18_n678));
   OAI2BB2XL U1099 (.Y(n1414), 
	.B1(FE_OFN16_n678), 
	.B0(n565), 
	.A1N(key_mem[873]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U1100 (.Y(n1413), 
	.B1(n678), 
	.B0(FE_PHN608_n564), 
	.A1N(FE_PHN3421_key_mem_874_), 
	.A0N(n678));
   OAI2BB2XL U1101 (.Y(n1412), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN615_n563), 
	.A1N(key_mem[875]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1102 (.Y(n1411), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN618_n562), 
	.A1N(key_mem[876]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1103 (.Y(n1410), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN621_n561), 
	.A1N(key_mem[877]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1104 (.Y(n1409), 
	.B1(FE_OFN16_n678), 
	.B0(n560), 
	.A1N(key_mem[878]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U1105 (.Y(n1408), 
	.B1(FE_OFN16_n678), 
	.B0(n559), 
	.A1N(FE_PHN3236_key_mem_879_), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U1106 (.Y(n1407), 
	.B1(FE_OFN16_n678), 
	.B0(n558), 
	.A1N(key_mem[880]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U1107 (.Y(n1406), 
	.B1(FE_OFN16_n678), 
	.B0(n557), 
	.A1N(key_mem[881]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U1108 (.Y(n1405), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN614_n556), 
	.A1N(key_mem[882]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1109 (.Y(n1404), 
	.B1(FE_OFN15_n678), 
	.B0(FE_PHN619_n555), 
	.A1N(key_mem[883]), 
	.A0N(FE_OFN15_n678));
   OAI2BB2XL U1110 (.Y(n1403), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN620_n554), 
	.A1N(key_mem[884]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U1111 (.Y(n1402), 
	.B1(FE_OFN17_n678), 
	.B0(FE_PHN616_n553), 
	.A1N(key_mem[885]), 
	.A0N(FE_OFN17_n678));
   OAI2BB2XL U1112 (.Y(n1401), 
	.B1(FE_OFN16_n678), 
	.B0(n552), 
	.A1N(key_mem[886]), 
	.A0N(FE_OFN16_n678));
   OAI2BB2XL U1113 (.Y(n1400), 
	.B1(FE_OFN16_n678), 
	.B0(FE_PHN624_n551), 
	.A1N(key_mem[887]), 
	.A0N(FE_OFN16_n678));
   AND3X2 U1114 (.Y(n686), 
	.C(FE_PHN116_round_ctr_reg_3_), 
	.B(n2873), 
	.A(n679));
   OAI2BB2XL U1115 (.Y(n2261), 
	.B1(FE_OFN12_n688), 
	.B0(FE_PHN401_n639), 
	.A1N(FE_PHN3085_key_mem_31_), 
	.A0N(FE_OFN12_n688));
   OAI2BB2XL U1116 (.Y(n2229), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN423_n607), 
	.A1N(key_mem[63]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1117 (.Y(n2197), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN342_n575), 
	.A1N(FE_PHN3201_key_mem_95_), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1118 (.Y(n2165), 
	.B1(FE_OFN12_n688), 
	.B0(FE_PHN622_n543), 
	.A1N(FE_PHN3208_key_mem_127_), 
	.A0N(FE_OFN12_n688));
   OAI2BB2XL U1119 (.Y(n2268), 
	.B1(FE_OFN12_n688), 
	.B0(FE_PHN406_n646), 
	.A1N(key_mem[24]), 
	.A0N(FE_OFN12_n688));
   OAI2BB2XL U1120 (.Y(n2236), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN404_n614), 
	.A1N(key_mem[56]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1121 (.Y(n2204), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN347_n582), 
	.A1N(key_mem[88]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1122 (.Y(n2172), 
	.B1(n688), 
	.B0(FE_PHN568_n550), 
	.A1N(key_mem[120]), 
	.A0N(n688));
   OAI2BB2XL U1123 (.Y(n2262), 
	.B1(FE_OFN12_n688), 
	.B0(FE_PHN408_n640), 
	.A1N(key_mem[30]), 
	.A0N(FE_OFN12_n688));
   OAI2BB2XL U1124 (.Y(n2230), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN422_n608), 
	.A1N(key_mem[62]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1125 (.Y(n2198), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN344_n576), 
	.A1N(key_mem[94]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1126 (.Y(n2166), 
	.B1(FE_OFN12_n688), 
	.B0(FE_PHN623_n544), 
	.A1N(FE_PHN3089_key_mem_126_), 
	.A0N(FE_OFN12_n688));
   OAI2BB2XL U1127 (.Y(n2263), 
	.B1(n688), 
	.B0(FE_PHN400_n641), 
	.A1N(key_mem[29]), 
	.A0N(n688));
   OAI2BB2XL U1128 (.Y(n2231), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN393_n609), 
	.A1N(key_mem[61]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1129 (.Y(n2199), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN343_n577), 
	.A1N(key_mem[93]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1130 (.Y(n2167), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN551_n545), 
	.A1N(key_mem[125]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1131 (.Y(n2264), 
	.B1(n688), 
	.B0(FE_PHN397_n642), 
	.A1N(key_mem[28]), 
	.A0N(n688));
   OAI2BB2XL U1132 (.Y(n2232), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN392_n610), 
	.A1N(key_mem[60]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1133 (.Y(n2200), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN345_n578), 
	.A1N(key_mem[92]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1134 (.Y(n2168), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN548_n546), 
	.A1N(key_mem[124]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1135 (.Y(n2265), 
	.B1(n688), 
	.B0(FE_PHN399_n643), 
	.A1N(key_mem[27]), 
	.A0N(n688));
   OAI2BB2XL U1136 (.Y(n2233), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN386_n611), 
	.A1N(key_mem[59]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1137 (.Y(n2201), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN346_n579), 
	.A1N(key_mem[91]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1138 (.Y(n2169), 
	.B1(n688), 
	.B0(FE_PHN544_n547), 
	.A1N(key_mem[123]), 
	.A0N(n688));
   OAI2BB2XL U1139 (.Y(n2266), 
	.B1(n688), 
	.B0(FE_PHN395_n644), 
	.A1N(key_mem[26]), 
	.A0N(n688));
   OAI2BB2XL U1140 (.Y(n2234), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN326_n612), 
	.A1N(key_mem[58]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1141 (.Y(n2202), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN547_n580), 
	.A1N(key_mem[90]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1142 (.Y(n2170), 
	.B1(n688), 
	.B0(FE_PHN418_n548), 
	.A1N(key_mem[122]), 
	.A0N(n688));
   OAI2BB2XL U1143 (.Y(n2267), 
	.B1(n688), 
	.B0(FE_PHN407_n645), 
	.A1N(key_mem[25]), 
	.A0N(n688));
   OAI2BB2XL U1144 (.Y(n2235), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN405_n613), 
	.A1N(key_mem[57]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1145 (.Y(n2203), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN349_n581), 
	.A1N(key_mem[89]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1146 (.Y(n2171), 
	.B1(n688), 
	.B0(FE_PHN567_n549), 
	.A1N(key_mem[121]), 
	.A0N(n688));
   OAI2BB2XL U1147 (.Y(n2292), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN553_n670), 
	.A1N(key_mem[0]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1148 (.Y(n2291), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN537_n669), 
	.A1N(key_mem[1]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1149 (.Y(n2290), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN550_n668), 
	.A1N(FE_PHN3248_key_mem_2_), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1150 (.Y(n2289), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN563_n667), 
	.A1N(key_mem[3]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1151 (.Y(n2288), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN562_n666), 
	.A1N(key_mem[4]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1152 (.Y(n2287), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN566_n665), 
	.A1N(key_mem[5]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1153 (.Y(n2286), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN572_n664), 
	.A1N(key_mem[6]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1154 (.Y(n2285), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN324_n663), 
	.A1N(key_mem[7]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1155 (.Y(n2284), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN325_n662), 
	.A1N(key_mem[8]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1156 (.Y(n2283), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN323_n661), 
	.A1N(key_mem[9]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1157 (.Y(n2282), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN541_n660), 
	.A1N(FE_PHN3206_key_mem_10_), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1158 (.Y(n2281), 
	.B1(n688), 
	.B0(FE_PHN554_n659), 
	.A1N(key_mem[11]), 
	.A0N(n688));
   OAI2BB2XL U1159 (.Y(n2280), 
	.B1(n688), 
	.B0(FE_PHN560_n658), 
	.A1N(key_mem[12]), 
	.A0N(n688));
   OAI2BB2XL U1160 (.Y(n2279), 
	.B1(n688), 
	.B0(FE_PHN552_n657), 
	.A1N(key_mem[13]), 
	.A0N(n688));
   OAI2BB2XL U1161 (.Y(n2278), 
	.B1(FE_OFN12_n688), 
	.B0(FE_PHN571_n656), 
	.A1N(key_mem[14]), 
	.A0N(FE_OFN12_n688));
   OAI2BB2XL U1162 (.Y(n2277), 
	.B1(FE_OFN12_n688), 
	.B0(FE_PHN327_n655), 
	.A1N(FE_PHN3283_key_mem_15_), 
	.A0N(FE_OFN12_n688));
   OAI2BB2XL U1163 (.Y(n2276), 
	.B1(FE_OFN12_n688), 
	.B0(FE_PHN573_n654), 
	.A1N(key_mem[16]), 
	.A0N(FE_OFN12_n688));
   OAI2BB2XL U1164 (.Y(n2275), 
	.B1(FE_OFN12_n688), 
	.B0(FE_PHN570_n653), 
	.A1N(key_mem[17]), 
	.A0N(FE_OFN12_n688));
   OAI2BB2XL U1165 (.Y(n2274), 
	.B1(FE_OFN12_n688), 
	.B0(FE_PHN558_n652), 
	.A1N(FE_PHN3194_key_mem_18_), 
	.A0N(FE_OFN12_n688));
   OAI2BB2XL U1166 (.Y(n2273), 
	.B1(FE_OFN12_n688), 
	.B0(FE_PHN569_n651), 
	.A1N(FE_PHN3188_key_mem_19_), 
	.A0N(FE_OFN12_n688));
   OAI2BB2XL U1167 (.Y(n2272), 
	.B1(FE_OFN12_n688), 
	.B0(FE_PHN579_n650), 
	.A1N(key_mem[20]), 
	.A0N(FE_OFN12_n688));
   OAI2BB2XL U1168 (.Y(n2271), 
	.B1(FE_OFN12_n688), 
	.B0(FE_PHN625_n649), 
	.A1N(key_mem[21]), 
	.A0N(FE_OFN12_n688));
   OAI2BB2XL U1169 (.Y(n2270), 
	.B1(FE_OFN12_n688), 
	.B0(FE_PHN564_n648), 
	.A1N(key_mem[22]), 
	.A0N(FE_OFN12_n688));
   OAI2BB2XL U1170 (.Y(n2269), 
	.B1(FE_OFN12_n688), 
	.B0(FE_PHN348_n647), 
	.A1N(key_mem[23]), 
	.A0N(FE_OFN12_n688));
   OAI2BB2XL U1171 (.Y(n2260), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN383_n638), 
	.A1N(key_mem[32]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1172 (.Y(n2259), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN380_n637), 
	.A1N(key_mem[33]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1173 (.Y(n2258), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN381_n636), 
	.A1N(key_mem[34]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1174 (.Y(n2257), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN379_n635), 
	.A1N(key_mem[35]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1175 (.Y(n2256), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN394_n634), 
	.A1N(key_mem[36]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1176 (.Y(n2255), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN391_n633), 
	.A1N(key_mem[37]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1177 (.Y(n2254), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN396_n632), 
	.A1N(key_mem[38]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1178 (.Y(n2253), 
	.B1(FE_OFN13_n688), 
	.B0(n631), 
	.A1N(key_mem[39]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1179 (.Y(n2252), 
	.B1(FE_OFN13_n688), 
	.B0(n630), 
	.A1N(key_mem[40]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1180 (.Y(n2251), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN705_n629), 
	.A1N(key_mem[41]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1181 (.Y(n2250), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN390_n628), 
	.A1N(key_mem[42]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1182 (.Y(n2249), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN398_n627), 
	.A1N(key_mem[43]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1183 (.Y(n2248), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN388_n626), 
	.A1N(key_mem[44]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1184 (.Y(n2247), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN387_n625), 
	.A1N(key_mem[45]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1185 (.Y(n2246), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN409_n624), 
	.A1N(key_mem[46]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1186 (.Y(n2245), 
	.B1(FE_OFN13_n688), 
	.B0(n623), 
	.A1N(key_mem[47]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1187 (.Y(n2244), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN403_n622), 
	.A1N(key_mem[48]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1188 (.Y(n2243), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN402_n621), 
	.A1N(key_mem[49]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1189 (.Y(n2242), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN384_n620), 
	.A1N(key_mem[50]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1190 (.Y(n2241), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN382_n619), 
	.A1N(key_mem[51]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1191 (.Y(n2240), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN389_n618), 
	.A1N(key_mem[52]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1192 (.Y(n2239), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN385_n617), 
	.A1N(key_mem[53]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1193 (.Y(n2238), 
	.B1(FE_OFN11_n688), 
	.B0(n616), 
	.A1N(key_mem[54]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1194 (.Y(n2237), 
	.B1(FE_OFN11_n688), 
	.B0(n615), 
	.A1N(key_mem[55]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1195 (.Y(n2228), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN540_n606), 
	.A1N(key_mem[64]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1196 (.Y(n2227), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN555_n605), 
	.A1N(key_mem[65]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1197 (.Y(n2226), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN538_n604), 
	.A1N(key_mem[66]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1198 (.Y(n2225), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN546_n603), 
	.A1N(key_mem[67]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1199 (.Y(n2224), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN557_n602), 
	.A1N(key_mem[68]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1200 (.Y(n2223), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN561_n601), 
	.A1N(key_mem[69]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1201 (.Y(n2222), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN578_n600), 
	.A1N(key_mem[70]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1202 (.Y(n2221), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN545_n599), 
	.A1N(key_mem[71]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1203 (.Y(n2220), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN559_n598), 
	.A1N(key_mem[72]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1204 (.Y(n2219), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN416_n597), 
	.A1N(FE_PHN3189_key_mem_73_), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1205 (.Y(n2218), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN565_n596), 
	.A1N(key_mem[74]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1206 (.Y(n2217), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN556_n595), 
	.A1N(key_mem[75]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1207 (.Y(n2216), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN575_n594), 
	.A1N(key_mem[76]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1208 (.Y(n2215), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN577_n593), 
	.A1N(key_mem[77]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1209 (.Y(n2214), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN420_n592), 
	.A1N(key_mem[78]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1210 (.Y(n2213), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN417_n591), 
	.A1N(key_mem[79]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1211 (.Y(n2212), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN421_n590), 
	.A1N(key_mem[80]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1212 (.Y(n2211), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN419_n589), 
	.A1N(key_mem[81]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1213 (.Y(n2210), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN543_n588), 
	.A1N(key_mem[82]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1214 (.Y(n2209), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN549_n587), 
	.A1N(key_mem[83]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1215 (.Y(n2208), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN542_n586), 
	.A1N(key_mem[84]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1216 (.Y(n2207), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN539_n585), 
	.A1N(key_mem[85]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1217 (.Y(n2206), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN576_n584), 
	.A1N(key_mem[86]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1218 (.Y(n2205), 
	.B1(n688), 
	.B0(FE_PHN574_n583), 
	.A1N(key_mem[87]), 
	.A0N(n688));
   OAI2BB2XL U1219 (.Y(n2196), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN609_n574), 
	.A1N(key_mem[96]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1220 (.Y(n2195), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN610_n573), 
	.A1N(key_mem[97]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1221 (.Y(n2194), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN612_n572), 
	.A1N(key_mem[98]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1222 (.Y(n2193), 
	.B1(FE_OFN13_n688), 
	.B0(FE_PHN606_n571), 
	.A1N(key_mem[99]), 
	.A0N(FE_OFN13_n688));
   OAI2BB2XL U1223 (.Y(n2192), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN617_n570), 
	.A1N(key_mem[100]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1224 (.Y(n2191), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN613_n569), 
	.A1N(key_mem[101]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1225 (.Y(n2190), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN605_n568), 
	.A1N(key_mem[102]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1226 (.Y(n2189), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN611_n567), 
	.A1N(key_mem[103]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1227 (.Y(n2188), 
	.B1(FE_OFN14_n688), 
	.B0(FE_PHN607_n566), 
	.A1N(key_mem[104]), 
	.A0N(FE_OFN14_n688));
   OAI2BB2XL U1228 (.Y(n2187), 
	.B1(n688), 
	.B0(n565), 
	.A1N(key_mem[105]), 
	.A0N(n688));
   OAI2BB2XL U1229 (.Y(n2186), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN608_n564), 
	.A1N(FE_PHN3185_key_mem_106_), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1230 (.Y(n2185), 
	.B1(n688), 
	.B0(FE_PHN615_n563), 
	.A1N(key_mem[107]), 
	.A0N(n688));
   OAI2BB2XL U1231 (.Y(n2184), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN618_n562), 
	.A1N(key_mem[108]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1232 (.Y(n2183), 
	.B1(n688), 
	.B0(FE_PHN621_n561), 
	.A1N(key_mem[109]), 
	.A0N(n688));
   OAI2BB2XL U1233 (.Y(n2182), 
	.B1(FE_OFN12_n688), 
	.B0(n560), 
	.A1N(key_mem[110]), 
	.A0N(FE_OFN12_n688));
   OAI2BB2XL U1234 (.Y(n2181), 
	.B1(FE_OFN12_n688), 
	.B0(n559), 
	.A1N(FE_PHN3187_key_mem_111_), 
	.A0N(FE_OFN12_n688));
   OAI2BB2XL U1235 (.Y(n2180), 
	.B1(FE_OFN12_n688), 
	.B0(n558), 
	.A1N(key_mem[112]), 
	.A0N(FE_OFN12_n688));
   OAI2BB2XL U1236 (.Y(n2179), 
	.B1(n688), 
	.B0(n557), 
	.A1N(key_mem[113]), 
	.A0N(n688));
   OAI2BB2XL U1237 (.Y(n2178), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN614_n556), 
	.A1N(key_mem[114]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1238 (.Y(n2177), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN619_n555), 
	.A1N(key_mem[115]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1239 (.Y(n2176), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN620_n554), 
	.A1N(key_mem[116]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1240 (.Y(n2175), 
	.B1(FE_OFN11_n688), 
	.B0(FE_PHN616_n553), 
	.A1N(key_mem[117]), 
	.A0N(FE_OFN11_n688));
   OAI2BB2XL U1241 (.Y(n2174), 
	.B1(FE_OFN12_n688), 
	.B0(n552), 
	.A1N(key_mem[118]), 
	.A0N(FE_OFN12_n688));
   OAI2BB2XL U1242 (.Y(n2173), 
	.B1(FE_OFN12_n688), 
	.B0(FE_PHN624_n551), 
	.A1N(key_mem[119]), 
	.A0N(FE_OFN12_n688));
   NOR3XL U1243 (.Y(n680), 
	.C(n2873), 
	.B(FE_PHN116_round_ctr_reg_3_), 
	.A(FE_PHN198_round_ctr_reg_0_));
   INVX1 U1244 (.Y(n2873), 
	.A(FE_PHN178_round_ctr_reg_2_));
   INVX1 U1245 (.Y(n2874), 
	.A(FE_PHN116_round_ctr_reg_3_));
   OAI2BB2XL U1246 (.Y(n2389), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN401_n639), 
	.A1N(sboxw[31]), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1247 (.Y(n2357), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN423_n607), 
	.A1N(FE_PHN743_prev_key1_reg_63_), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1248 (.Y(n2325), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN342_n575), 
	.A1N(FE_PHN940_prev_key1_reg_95_), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1249 (.Y(n2293), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN622_n543), 
	.A1N(FE_PHN1434_prev_key1_reg_127_), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1250 (.Y(n2396), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN406_n646), 
	.A1N(sboxw[24]), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1251 (.Y(n2364), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN404_n614), 
	.A1N(prev_key1_reg[56]), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1252 (.Y(n2332), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN347_n582), 
	.A1N(FE_PHN979_prev_key1_reg_88_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1253 (.Y(n2300), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN568_n550), 
	.A1N(FE_PHN1416_prev_key1_reg_120_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1254 (.Y(n2390), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN408_n640), 
	.A1N(sboxw[30]), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1255 (.Y(n2358), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN422_n608), 
	.A1N(FE_PHN740_prev_key1_reg_62_), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1256 (.Y(n2326), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN344_n576), 
	.A1N(FE_PHN933_prev_key1_reg_94_), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1257 (.Y(n2294), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN623_n544), 
	.A1N(prev_key1_reg[126]), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1258 (.Y(n2391), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN400_n641), 
	.A1N(sboxw[29]), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1259 (.Y(n2359), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN393_n609), 
	.A1N(FE_PHN896_prev_key1_reg_61_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1260 (.Y(n2327), 
	.B1(n683), 
	.B0(FE_PHN343_n577), 
	.A1N(FE_PHN757_prev_key1_reg_93_), 
	.A0N(n683));
   OAI2BB2XL U1261 (.Y(n2295), 
	.B1(n683), 
	.B0(FE_PHN551_n545), 
	.A1N(FE_PHN1391_prev_key1_reg_125_), 
	.A0N(n683));
   OAI2BB2XL U1262 (.Y(n2392), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN397_n642), 
	.A1N(sboxw[28]), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1263 (.Y(n2360), 
	.B1(n683), 
	.B0(FE_PHN392_n610), 
	.A1N(FE_PHN741_prev_key1_reg_60_), 
	.A0N(n683));
   OAI2BB2XL U1264 (.Y(n2328), 
	.B1(n683), 
	.B0(FE_PHN345_n578), 
	.A1N(FE_PHN919_prev_key1_reg_92_), 
	.A0N(n683));
   OAI2BB2XL U1265 (.Y(n2296), 
	.B1(n683), 
	.B0(FE_PHN548_n546), 
	.A1N(FE_PHN1421_prev_key1_reg_124_), 
	.A0N(n683));
   OAI2BB2XL U1266 (.Y(n2393), 
	.B1(n683), 
	.B0(FE_PHN399_n643), 
	.A1N(sboxw[27]), 
	.A0N(n683));
   OAI2BB2XL U1267 (.Y(n2361), 
	.B1(n683), 
	.B0(FE_PHN386_n611), 
	.A1N(FE_PHN745_prev_key1_reg_59_), 
	.A0N(n683));
   OAI2BB2XL U1268 (.Y(n2329), 
	.B1(n683), 
	.B0(FE_PHN346_n579), 
	.A1N(FE_PHN921_prev_key1_reg_91_), 
	.A0N(n683));
   OAI2BB2XL U1269 (.Y(n2297), 
	.B1(n683), 
	.B0(FE_PHN544_n547), 
	.A1N(FE_PHN1413_prev_key1_reg_123_), 
	.A0N(n683));
   OAI2BB2XL U1270 (.Y(n2394), 
	.B1(n683), 
	.B0(FE_PHN395_n644), 
	.A1N(sboxw[26]), 
	.A0N(n683));
   OAI2BB2XL U1271 (.Y(n2362), 
	.B1(n683), 
	.B0(FE_PHN326_n612), 
	.A1N(FE_PHN746_prev_key1_reg_58_), 
	.A0N(n683));
   OAI2BB2XL U1272 (.Y(n2330), 
	.B1(n683), 
	.B0(FE_PHN547_n580), 
	.A1N(FE_PHN924_prev_key1_reg_90_), 
	.A0N(n683));
   OAI2BB2XL U1273 (.Y(n2298), 
	.B1(n683), 
	.B0(FE_PHN418_n548), 
	.A1N(FE_PHN1392_prev_key1_reg_122_), 
	.A0N(n683));
   OAI2BB2XL U1274 (.Y(n2395), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN407_n645), 
	.A1N(sboxw[25]), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1275 (.Y(n2363), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN405_n613), 
	.A1N(FE_PHN744_prev_key1_reg_57_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1276 (.Y(n2331), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN349_n581), 
	.A1N(FE_PHN922_prev_key1_reg_89_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1277 (.Y(n2299), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN567_n549), 
	.A1N(FE_PHN1395_prev_key1_reg_121_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1278 (.Y(n2420), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN553_n670), 
	.A1N(FE_PHN1959_keymem_sboxw_0_), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1279 (.Y(n2419), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN537_n669), 
	.A1N(sboxw[1]), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1280 (.Y(n2418), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN550_n668), 
	.A1N(sboxw[2]), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1281 (.Y(n2417), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN563_n667), 
	.A1N(sboxw[3]), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1282 (.Y(n2416), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN562_n666), 
	.A1N(FE_PHN2003_keymem_sboxw_4_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1283 (.Y(n2415), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN566_n665), 
	.A1N(FE_PHN2006_keymem_sboxw_5_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1284 (.Y(n2414), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN572_n664), 
	.A1N(sboxw[6]), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1285 (.Y(n2413), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN324_n663), 
	.A1N(sboxw[7]), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1286 (.Y(n2412), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN325_n662), 
	.A1N(FE_PHN2001_keymem_sboxw_8_), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1287 (.Y(n2411), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN323_n661), 
	.A1N(sboxw[9]), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1288 (.Y(n2410), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN541_n660), 
	.A1N(FE_PHN1962_keymem_sboxw_10_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1289 (.Y(n2409), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN554_n659), 
	.A1N(sboxw[11]), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1290 (.Y(n2408), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN560_n658), 
	.A1N(FE_PHN2004_keymem_sboxw_12_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1291 (.Y(n2407), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN552_n657), 
	.A1N(sboxw[13]), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1292 (.Y(n2406), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN571_n656), 
	.A1N(sboxw[14]), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1293 (.Y(n2405), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN327_n655), 
	.A1N(sboxw[15]), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1294 (.Y(n2404), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN573_n654), 
	.A1N(sboxw[16]), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1295 (.Y(n2403), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN570_n653), 
	.A1N(FE_PHN1998_keymem_sboxw_17_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1296 (.Y(n2402), 
	.B1(n683), 
	.B0(FE_PHN558_n652), 
	.A1N(FE_PHN1958_keymem_sboxw_18_), 
	.A0N(n683));
   OAI2BB2XL U1297 (.Y(n2401), 
	.B1(n683), 
	.B0(FE_PHN569_n651), 
	.A1N(sboxw[19]), 
	.A0N(n683));
   OAI2BB2XL U1298 (.Y(n2400), 
	.B1(n683), 
	.B0(FE_PHN579_n650), 
	.A1N(FE_PHN2005_keymem_sboxw_20_), 
	.A0N(n683));
   OAI2BB2XL U1299 (.Y(n2399), 
	.B1(n683), 
	.B0(FE_PHN625_n649), 
	.A1N(sboxw[21]), 
	.A0N(n683));
   OAI2BB2XL U1300 (.Y(n2398), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN564_n648), 
	.A1N(FE_PHN1965_keymem_sboxw_22_), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1301 (.Y(n2397), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN348_n647), 
	.A1N(sboxw[23]), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1303 (.Y(n2388), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN383_n638), 
	.A1N(FE_PHN1079_prev_key1_reg_32_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1304 (.Y(n2387), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN380_n637), 
	.A1N(FE_PHN1060_prev_key1_reg_33_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1305 (.Y(n2386), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN381_n636), 
	.A1N(FE_PHN1044_prev_key1_reg_34_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1306 (.Y(n2385), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN379_n635), 
	.A1N(FE_PHN1063_prev_key1_reg_35_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1307 (.Y(n2384), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN394_n634), 
	.A1N(FE_PHN1053_prev_key1_reg_36_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1308 (.Y(n2383), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN391_n633), 
	.A1N(FE_PHN1056_prev_key1_reg_37_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1309 (.Y(n2382), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN396_n632), 
	.A1N(FE_PHN1055_prev_key1_reg_38_), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1310 (.Y(n2381), 
	.B1(FE_OFN33_n683), 
	.B0(n631), 
	.A1N(FE_PHN1049_prev_key1_reg_39_), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1311 (.Y(n2380), 
	.B1(FE_OFN32_n683), 
	.B0(n630), 
	.A1N(FE_PHN1051_prev_key1_reg_40_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1312 (.Y(n2379), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN705_n629), 
	.A1N(FE_PHN1058_prev_key1_reg_41_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1313 (.Y(n2378), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN390_n628), 
	.A1N(FE_PHN1054_prev_key1_reg_42_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1314 (.Y(n2377), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN398_n627), 
	.A1N(FE_PHN1048_prev_key1_reg_43_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1315 (.Y(n2376), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN388_n626), 
	.A1N(FE_PHN1087_prev_key1_reg_44_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1316 (.Y(n2375), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN387_n625), 
	.A1N(FE_PHN1064_prev_key1_reg_45_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1317 (.Y(n2374), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN409_n624), 
	.A1N(prev_key1_reg[46]), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1318 (.Y(n2373), 
	.B1(FE_OFN33_n683), 
	.B0(n623), 
	.A1N(FE_PHN1062_prev_key1_reg_47_), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1319 (.Y(n2372), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN403_n622), 
	.A1N(prev_key1_reg[48]), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1320 (.Y(n2371), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN402_n621), 
	.A1N(FE_PHN1067_prev_key1_reg_49_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1321 (.Y(n2370), 
	.B1(n683), 
	.B0(FE_PHN384_n620), 
	.A1N(FE_PHN1074_prev_key1_reg_50_), 
	.A0N(n683));
   OAI2BB2XL U1322 (.Y(n2369), 
	.B1(n683), 
	.B0(FE_PHN382_n619), 
	.A1N(FE_PHN1052_prev_key1_reg_51_), 
	.A0N(n683));
   OAI2BB2XL U1323 (.Y(n2368), 
	.B1(n683), 
	.B0(FE_PHN389_n618), 
	.A1N(FE_PHN1043_prev_key1_reg_52_), 
	.A0N(n683));
   OAI2BB2XL U1324 (.Y(n2367), 
	.B1(n683), 
	.B0(FE_PHN385_n617), 
	.A1N(FE_PHN1230_prev_key1_reg_53_), 
	.A0N(n683));
   OAI2BB2XL U1325 (.Y(n2366), 
	.B1(FE_OFN31_n683), 
	.B0(n616), 
	.A1N(FE_PHN1050_prev_key1_reg_54_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1326 (.Y(n2365), 
	.B1(FE_OFN31_n683), 
	.B0(n615), 
	.A1N(FE_PHN1057_prev_key1_reg_55_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1327 (.Y(n2356), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN540_n606), 
	.A1N(FE_PHN1441_prev_key1_reg_64_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1328 (.Y(n2355), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN555_n605), 
	.A1N(FE_PHN1394_prev_key1_reg_65_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1329 (.Y(n2354), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN538_n604), 
	.A1N(FE_PHN1442_prev_key1_reg_66_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1330 (.Y(n2353), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN546_n603), 
	.A1N(FE_PHN1444_prev_key1_reg_67_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1331 (.Y(n2352), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN557_n602), 
	.A1N(FE_PHN1446_prev_key1_reg_68_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1332 (.Y(n2351), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN561_n601), 
	.A1N(FE_PHN1445_prev_key1_reg_69_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1333 (.Y(n2350), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN578_n600), 
	.A1N(prev_key1_reg[70]), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1334 (.Y(n2349), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN545_n599), 
	.A1N(FE_PHN1406_prev_key1_reg_71_), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1335 (.Y(n2348), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN559_n598), 
	.A1N(FE_PHN1404_prev_key1_reg_72_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1336 (.Y(n2347), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN416_n597), 
	.A1N(FE_PHN1401_prev_key1_reg_73_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1337 (.Y(n2346), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN565_n596), 
	.A1N(FE_PHN1408_prev_key1_reg_74_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1338 (.Y(n2345), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN556_n595), 
	.A1N(FE_PHN1415_prev_key1_reg_75_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1339 (.Y(n2344), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN575_n594), 
	.A1N(FE_PHN1429_prev_key1_reg_76_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1340 (.Y(n2343), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN577_n593), 
	.A1N(FE_PHN1397_prev_key1_reg_77_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1341 (.Y(n2342), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN420_n592), 
	.A1N(FE_PHN1402_prev_key1_reg_78_), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1342 (.Y(n2341), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN417_n591), 
	.A1N(FE_PHN1393_prev_key1_reg_79_), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1343 (.Y(n2340), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN421_n590), 
	.A1N(FE_PHN1414_prev_key1_reg_80_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1344 (.Y(n2339), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN419_n589), 
	.A1N(FE_PHN1425_prev_key1_reg_81_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1345 (.Y(n2338), 
	.B1(n683), 
	.B0(FE_PHN543_n588), 
	.A1N(FE_PHN1405_prev_key1_reg_82_), 
	.A0N(n683));
   OAI2BB2XL U1346 (.Y(n2337), 
	.B1(n683), 
	.B0(FE_PHN549_n587), 
	.A1N(FE_PHN1388_prev_key1_reg_83_), 
	.A0N(n683));
   OAI2BB2XL U1347 (.Y(n2336), 
	.B1(n683), 
	.B0(FE_PHN542_n586), 
	.A1N(FE_PHN1375_prev_key1_reg_84_), 
	.A0N(n683));
   OAI2BB2XL U1348 (.Y(n2335), 
	.B1(n683), 
	.B0(FE_PHN539_n585), 
	.A1N(FE_PHN1412_prev_key1_reg_85_), 
	.A0N(n683));
   OAI2BB2XL U1349 (.Y(n2334), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN576_n584), 
	.A1N(FE_PHN360_prev_key1_reg_86_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1350 (.Y(n2333), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN574_n583), 
	.A1N(FE_PHN359_prev_key1_reg_87_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1351 (.Y(n2324), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN609_n574), 
	.A1N(FE_PHN1231_prev_key1_reg_96_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1352 (.Y(n2323), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN610_n573), 
	.A1N(FE_PHN1239_prev_key1_reg_97_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1353 (.Y(n2322), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN612_n572), 
	.A1N(FE_PHN1238_prev_key1_reg_98_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1354 (.Y(n2321), 
	.B1(FE_OFN32_n683), 
	.B0(FE_PHN606_n571), 
	.A1N(FE_PHN1245_prev_key1_reg_99_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1355 (.Y(n2320), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN617_n570), 
	.A1N(FE_PHN1225_prev_key1_reg_100_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1356 (.Y(n2319), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN613_n569), 
	.A1N(FE_PHN1229_prev_key1_reg_101_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1357 (.Y(n2318), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN605_n568), 
	.A1N(FE_PHN1220_prev_key1_reg_102_), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1358 (.Y(n2317), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN611_n567), 
	.A1N(FE_PHN1224_prev_key1_reg_103_), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1359 (.Y(n2316), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN607_n566), 
	.A1N(FE_PHN1223_prev_key1_reg_104_), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1360 (.Y(n2315), 
	.B1(FE_OFN32_n683), 
	.B0(n565), 
	.A1N(FE_PHN1252_prev_key1_reg_105_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1361 (.Y(n2314), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN608_n564), 
	.A1N(FE_PHN1233_prev_key1_reg_106_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1362 (.Y(n2313), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN615_n563), 
	.A1N(FE_PHN1232_prev_key1_reg_107_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1363 (.Y(n2312), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN618_n562), 
	.A1N(FE_PHN1251_prev_key1_reg_108_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1364 (.Y(n2311), 
	.B1(FE_OFN31_n683), 
	.B0(FE_PHN621_n561), 
	.A1N(FE_PHN1234_prev_key1_reg_109_), 
	.A0N(FE_OFN31_n683));
   OAI2BB2XL U1365 (.Y(n2310), 
	.B1(FE_OFN33_n683), 
	.B0(n560), 
	.A1N(FE_PHN1219_prev_key1_reg_110_), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1366 (.Y(n2309), 
	.B1(FE_OFN33_n683), 
	.B0(n559), 
	.A1N(FE_PHN1221_prev_key1_reg_111_), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1367 (.Y(n2308), 
	.B1(FE_OFN32_n683), 
	.B0(n558), 
	.A1N(FE_PHN1256_prev_key1_reg_112_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1368 (.Y(n2307), 
	.B1(FE_OFN32_n683), 
	.B0(n557), 
	.A1N(FE_PHN1236_prev_key1_reg_113_), 
	.A0N(FE_OFN32_n683));
   OAI2BB2XL U1369 (.Y(n2306), 
	.B1(n683), 
	.B0(FE_PHN614_n556), 
	.A1N(FE_PHN1226_prev_key1_reg_114_), 
	.A0N(n683));
   OAI2BB2XL U1370 (.Y(n2305), 
	.B1(n683), 
	.B0(FE_PHN619_n555), 
	.A1N(FE_PHN1244_prev_key1_reg_115_), 
	.A0N(n683));
   OAI2BB2XL U1371 (.Y(n2304), 
	.B1(n683), 
	.B0(FE_PHN620_n554), 
	.A1N(FE_PHN1249_prev_key1_reg_116_), 
	.A0N(n683));
   OAI2BB2XL U1372 (.Y(n2303), 
	.B1(n683), 
	.B0(FE_PHN616_n553), 
	.A1N(FE_PHN1235_prev_key1_reg_117_), 
	.A0N(n683));
   OAI2BB2XL U1373 (.Y(n2302), 
	.B1(FE_OFN33_n683), 
	.B0(n552), 
	.A1N(FE_PHN1313_prev_key1_reg_118_), 
	.A0N(FE_OFN33_n683));
   OAI2BB2XL U1374 (.Y(n2301), 
	.B1(FE_OFN33_n683), 
	.B0(FE_PHN624_n551), 
	.A1N(FE_PHN1314_prev_key1_reg_119_), 
	.A0N(FE_OFN33_n683));
   NAND3XL U1375 (.Y(n677), 
	.C(FE_PHN112_round_ctr_reg_1_), 
	.B(n2874), 
	.A(FE_PHN198_round_ctr_reg_0_));
   NAND4X1 U1376 (.Y(n689), 
	.D(n2873), 
	.C(FE_PHN411_n6), 
	.B(FE_PHN112_round_ctr_reg_1_), 
	.A(FE_PHN116_round_ctr_reg_3_));
   XOR2X1 U1377 (.Y(n720), 
	.B(new_sboxw[2]), 
	.A(FE_PHN1233_prev_key1_reg_106_));
   XOR2X1 U1378 (.Y(n717), 
	.B(new_sboxw[5]), 
	.A(FE_PHN1234_prev_key1_reg_109_));
   XOR2X1 U1379 (.Y(n715), 
	.B(new_sboxw[7]), 
	.A(FE_PHN1221_prev_key1_reg_111_));
   XOR2X1 U1380 (.Y(n728), 
	.B(new_sboxw[26]), 
	.A(FE_PHN1238_prev_key1_reg_98_));
   XOR2X1 U1381 (.Y(n722), 
	.B(new_sboxw[0]), 
	.A(FE_PHN1223_prev_key1_reg_104_));
   XOR2X1 U1382 (.Y(n721), 
	.B(new_sboxw[1]), 
	.A(FE_PHN1252_prev_key1_reg_105_));
   XOR2X1 U1383 (.Y(n719), 
	.B(new_sboxw[3]), 
	.A(FE_PHN1232_prev_key1_reg_107_));
   XOR2X1 U1384 (.Y(n718), 
	.B(new_sboxw[4]), 
	.A(FE_PHN1251_prev_key1_reg_108_));
   XOR2X1 U1385 (.Y(n730), 
	.B(new_sboxw[24]), 
	.A(FE_PHN1231_prev_key1_reg_96_));
   XOR2X1 U1386 (.Y(n729), 
	.B(new_sboxw[25]), 
	.A(FE_PHN1239_prev_key1_reg_97_));
   XOR2X1 U1387 (.Y(n727), 
	.B(new_sboxw[27]), 
	.A(FE_PHN1245_prev_key1_reg_99_));
   XOR2X1 U1388 (.Y(n692), 
	.B(new_sboxw[23]), 
	.A(FE_PHN912_rcon_reg_7_));
   XOR2X1 U1389 (.Y(n696), 
	.B(new_sboxw[21]), 
	.A(FE_PHN1241_rcon_reg_5_));
   XOR2X1 U1390 (.Y(n702), 
	.B(new_sboxw[18]), 
	.A(FE_PHN1033_rcon_reg_2_));
   XOR2X1 U1391 (.Y(n706), 
	.B(new_sboxw[16]), 
	.A(FE_PHN1034_rcon_reg_0_));
   XOR2X1 U1392 (.Y(n700), 
	.B(new_sboxw[19]), 
	.A(FE_PHN1036_rcon_reg_3_));
   XOR2X1 U1393 (.Y(n704), 
	.B(new_sboxw[17]), 
	.A(FE_PHN1263_rcon_reg_1_));
   XOR2X1 U1394 (.Y(n698), 
	.B(new_sboxw[20]), 
	.A(FE_PHN1257_rcon_reg_4_));
   XNOR2X1 U1395 (.Y(n810), 
	.B(n730), 
	.A(n874));
   XNOR2X1 U1396 (.Y(n874), 
	.B(FE_PHN1441_prev_key1_reg_64_), 
	.A(FE_PHN1079_prev_key1_reg_32_));
   XNOR2X1 U1397 (.Y(n809), 
	.B(n729), 
	.A(n872));
   XNOR2X1 U1398 (.Y(n872), 
	.B(FE_PHN1394_prev_key1_reg_65_), 
	.A(FE_PHN1060_prev_key1_reg_33_));
   XNOR2X1 U1399 (.Y(n808), 
	.B(n728), 
	.A(n870));
   XNOR2X1 U1400 (.Y(n870), 
	.B(FE_PHN1442_prev_key1_reg_66_), 
	.A(FE_PHN1044_prev_key1_reg_34_));
   XNOR2X1 U1401 (.Y(n807), 
	.B(n727), 
	.A(n868));
   XNOR2X1 U1402 (.Y(n868), 
	.B(FE_PHN1444_prev_key1_reg_67_), 
	.A(FE_PHN1063_prev_key1_reg_35_));
   XNOR2X1 U1403 (.Y(n802), 
	.B(n722), 
	.A(n858));
   XNOR2X1 U1404 (.Y(n858), 
	.B(FE_PHN1404_prev_key1_reg_72_), 
	.A(FE_PHN1051_prev_key1_reg_40_));
   XNOR2X1 U1405 (.Y(n801), 
	.B(n721), 
	.A(n856));
   XNOR2X1 U1406 (.Y(n856), 
	.B(FE_PHN1401_prev_key1_reg_73_), 
	.A(FE_PHN1058_prev_key1_reg_41_));
   XNOR2X1 U1407 (.Y(n800), 
	.B(n720), 
	.A(n854));
   XNOR2X1 U1408 (.Y(n854), 
	.B(FE_PHN1408_prev_key1_reg_74_), 
	.A(FE_PHN1054_prev_key1_reg_42_));
   XNOR2X1 U1409 (.Y(n799), 
	.B(n719), 
	.A(n852));
   XNOR2X1 U1410 (.Y(n852), 
	.B(FE_PHN1415_prev_key1_reg_75_), 
	.A(FE_PHN1048_prev_key1_reg_43_));
   XNOR2X1 U1411 (.Y(n798), 
	.B(n718), 
	.A(n850));
   XNOR2X1 U1412 (.Y(n850), 
	.B(FE_PHN1429_prev_key1_reg_76_), 
	.A(FE_PHN1087_prev_key1_reg_44_));
   XNOR2X1 U1413 (.Y(n797), 
	.B(n717), 
	.A(n848));
   XNOR2X1 U1414 (.Y(n848), 
	.B(FE_PHN1397_prev_key1_reg_77_), 
	.A(FE_PHN1064_prev_key1_reg_45_));
   XNOR2X1 U1415 (.Y(n795), 
	.B(n715), 
	.A(n844));
   XNOR2X1 U1416 (.Y(n844), 
	.B(FE_PHN1393_prev_key1_reg_79_), 
	.A(FE_PHN1062_prev_key1_reg_47_));
   OAI2BB2X1 U1417 (.Y(n1370), 
	.B1(n676), 
	.B0(FE_PHN395_n644), 
	.A1N(key_mem[922]), 
	.A0N(n676));
   OAI2BB2X1 U1418 (.Y(n1242), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN395_n644), 
	.A1N(FE_PHN1772_key_mem_1050_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1419 (.Y(n1114), 
	.B1(n672), 
	.B0(FE_PHN395_n644), 
	.A1N(key_mem[1178]), 
	.A0N(n672));
   OAI2BB2X1 U1420 (.Y(n986), 
	.B1(n1), 
	.B0(FE_PHN395_n644), 
	.A1N(key_mem[1306]), 
	.A0N(n1));
   AOI22X1 U1422 (.Y(n580), 
	.B1(n2655), 
	.B0(key[90]), 
	.A1(n736), 
	.A0(FE_OFN90_n690));
   AOI22X1 U1424 (.Y(n639), 
	.B1(n2685), 
	.B0(key[31]), 
	.A1(n811), 
	.A0(FE_OFN91_n690));
   XNOR2X1 U1425 (.Y(n811), 
	.B(n731), 
	.A(n812));
   XNOR2X1 U1426 (.Y(n812), 
	.B(sboxw[31]), 
	.A(FE_PHN743_prev_key1_reg_63_));
   AOI22X1 U1428 (.Y(n607), 
	.B1(n2669), 
	.B0(key[63]), 
	.A1(n763), 
	.A0(FE_OFN91_n690));
   XNOR2X1 U1429 (.Y(n763), 
	.B(n765), 
	.A(n764));
   XNOR2X1 U1430 (.Y(n764), 
	.B(n692), 
	.A(FE_PHN743_prev_key1_reg_63_));
   AOI22X1 U1433 (.Y(n646), 
	.B1(n2688), 
	.B0(key[24]), 
	.A1(n825), 
	.A0(FE_OFN91_n690));
   XNOR2X1 U1434 (.Y(n825), 
	.B(n738), 
	.A(n826));
   XNOR2X1 U1435 (.Y(n826), 
	.B(sboxw[24]), 
	.A(prev_key1_reg[56]));
   AOI22X1 U1437 (.Y(n614), 
	.B1(n2672), 
	.B0(key[56]), 
	.A1(n784), 
	.A0(FE_OFN91_n690));
   XNOR2X1 U1438 (.Y(n784), 
	.B(n786), 
	.A(n785));
   XNOR2X1 U1439 (.Y(n785), 
	.B(n706), 
	.A(prev_key1_reg[56]));
   AOI22X1 U1441 (.Y(n641), 
	.B1(n2686), 
	.B0(key[29]), 
	.A1(n815), 
	.A0(FE_OFN90_n690));
   XNOR2X1 U1442 (.Y(n815), 
	.B(n733), 
	.A(n816));
   XNOR2X1 U1443 (.Y(n816), 
	.B(sboxw[29]), 
	.A(FE_PHN896_prev_key1_reg_61_));
   AOI22X1 U1445 (.Y(n609), 
	.B1(n2670), 
	.B0(key[61]), 
	.A1(n769), 
	.A0(FE_OFN90_n690));
   XNOR2X1 U1446 (.Y(n769), 
	.B(n771), 
	.A(n770));
   XNOR2X1 U1447 (.Y(n770), 
	.B(n696), 
	.A(FE_PHN896_prev_key1_reg_61_));
   AOI22X1 U1449 (.Y(n642), 
	.B1(n2686), 
	.B0(key[28]), 
	.A1(n817), 
	.A0(FE_OFN90_n690));
   XNOR2X1 U1450 (.Y(n817), 
	.B(n734), 
	.A(n818));
   XNOR2X1 U1451 (.Y(n818), 
	.B(sboxw[28]), 
	.A(FE_PHN741_prev_key1_reg_60_));
   AOI22X1 U1453 (.Y(n643), 
	.B1(n2687), 
	.B0(key[27]), 
	.A1(n819), 
	.A0(FE_OFN90_n690));
   XNOR2X1 U1454 (.Y(n819), 
	.B(n735), 
	.A(n820));
   XNOR2X1 U1455 (.Y(n820), 
	.B(sboxw[27]), 
	.A(FE_PHN745_prev_key1_reg_59_));
   AOI22X1 U1457 (.Y(n611), 
	.B1(n2671), 
	.B0(key[59]), 
	.A1(n775), 
	.A0(FE_OFN90_n690));
   XNOR2X1 U1458 (.Y(n775), 
	.B(n777), 
	.A(n776));
   XNOR2X1 U1459 (.Y(n776), 
	.B(n700), 
	.A(FE_PHN745_prev_key1_reg_59_));
   AOI22X1 U1461 (.Y(n644), 
	.B1(n2687), 
	.B0(key[26]), 
	.A1(n821), 
	.A0(FE_OFN90_n690));
   XNOR2X1 U1462 (.Y(n821), 
	.B(n736), 
	.A(n822));
   XNOR2X1 U1463 (.Y(n822), 
	.B(sboxw[26]), 
	.A(FE_PHN746_prev_key1_reg_58_));
   AOI22X1 U1465 (.Y(n612), 
	.B1(n2671), 
	.B0(key[58]), 
	.A1(n778), 
	.A0(FE_OFN90_n690));
   XNOR2X1 U1466 (.Y(n778), 
	.B(n780), 
	.A(n779));
   XNOR2X1 U1467 (.Y(n779), 
	.B(n702), 
	.A(FE_PHN746_prev_key1_reg_58_));
   AOI22X1 U1469 (.Y(n645), 
	.B1(n2688), 
	.B0(key[25]), 
	.A1(n823), 
	.A0(FE_OFN91_n690));
   XNOR2X1 U1470 (.Y(n823), 
	.B(n737), 
	.A(n824));
   XNOR2X1 U1471 (.Y(n824), 
	.B(sboxw[25]), 
	.A(FE_PHN744_prev_key1_reg_57_));
   AOI22X1 U1473 (.Y(n613), 
	.B1(n2672), 
	.B0(key[57]), 
	.A1(n781), 
	.A0(FE_OFN91_n690));
   XNOR2X1 U1474 (.Y(n781), 
	.B(n783), 
	.A(n782));
   XNOR2X1 U1475 (.Y(n782), 
	.B(n704), 
	.A(FE_PHN744_prev_key1_reg_57_));
   AOI22X1 U1477 (.Y(n670), 
	.B1(n2699), 
	.B0(key[0]), 
	.A1(n873), 
	.A0(FE_OFN91_n690));
   XOR2X1 U1478 (.Y(n873), 
	.B(n810), 
	.A(FE_PHN1959_keymem_sboxw_0_));
   AOI22X1 U1480 (.Y(n669), 
	.B1(n2699), 
	.B0(key[1]), 
	.A1(n871), 
	.A0(FE_OFN91_n690));
   XOR2X1 U1481 (.Y(n871), 
	.B(n809), 
	.A(sboxw[1]));
   AOI22X1 U1483 (.Y(n668), 
	.B1(n2699), 
	.B0(key[2]), 
	.A1(n869), 
	.A0(FE_OFN91_n690));
   XOR2X1 U1484 (.Y(n869), 
	.B(n808), 
	.A(sboxw[2]));
   AOI22X1 U1486 (.Y(n667), 
	.B1(n2699), 
	.B0(key[3]), 
	.A1(n867), 
	.A0(FE_OFN91_n690));
   XOR2X1 U1487 (.Y(n867), 
	.B(n807), 
	.A(sboxw[3]));
   AOI22X1 U1489 (.Y(n662), 
	.B1(n2696), 
	.B0(key[8]), 
	.A1(n857), 
	.A0(FE_OFN91_n690));
   XOR2X1 U1490 (.Y(n857), 
	.B(n802), 
	.A(FE_PHN2001_keymem_sboxw_8_));
   AOI22X1 U1492 (.Y(n661), 
	.B1(n2696), 
	.B0(key[9]), 
	.A1(n855), 
	.A0(FE_OFN91_n690));
   XOR2X1 U1493 (.Y(n855), 
	.B(n801), 
	.A(sboxw[9]));
   AOI22X1 U1495 (.Y(n660), 
	.B1(n2695), 
	.B0(key[10]), 
	.A1(n853), 
	.A0(FE_OFN90_n690));
   XOR2X1 U1496 (.Y(n853), 
	.B(n800), 
	.A(FE_PHN1962_keymem_sboxw_10_));
   AOI22X1 U1498 (.Y(n659), 
	.B1(n2695), 
	.B0(key[11]), 
	.A1(n851), 
	.A0(FE_OFN90_n690));
   XOR2X1 U1499 (.Y(n851), 
	.B(n799), 
	.A(sboxw[11]));
   AOI22X1 U1501 (.Y(n658), 
	.B1(n2694), 
	.B0(key[12]), 
	.A1(n849), 
	.A0(FE_OFN90_n690));
   XOR2X1 U1502 (.Y(n849), 
	.B(n798), 
	.A(FE_PHN2004_keymem_sboxw_12_));
   AOI22X1 U1504 (.Y(n657), 
	.B1(n2694), 
	.B0(key[13]), 
	.A1(n847), 
	.A0(FE_OFN90_n690));
   XOR2X1 U1505 (.Y(n847), 
	.B(n797), 
	.A(sboxw[13]));
   AOI22X1 U1507 (.Y(n655), 
	.B1(n2693), 
	.B0(key[15]), 
	.A1(n843), 
	.A0(FE_OFN91_n690));
   XOR2X1 U1508 (.Y(n843), 
	.B(n795), 
	.A(sboxw[15]));
   XOR2X1 U1509 (.Y(n712), 
	.B(new_sboxw[10]), 
	.A(FE_PHN1226_prev_key1_reg_114_));
   XOR2X1 U1510 (.Y(n709), 
	.B(new_sboxw[13]), 
	.A(FE_PHN1235_prev_key1_reg_117_));
   XOR2X1 U1511 (.Y(n707), 
	.B(new_sboxw[15]), 
	.A(FE_PHN1314_prev_key1_reg_119_));
   XOR2X1 U1512 (.Y(n725), 
	.B(new_sboxw[29]), 
	.A(FE_PHN1229_prev_key1_reg_101_));
   XOR2X1 U1513 (.Y(n723), 
	.B(new_sboxw[31]), 
	.A(FE_PHN1224_prev_key1_reg_103_));
   XOR2X1 U1514 (.Y(n716), 
	.B(new_sboxw[6]), 
	.A(FE_PHN1219_prev_key1_reg_110_));
   XOR2X1 U1515 (.Y(n714), 
	.B(new_sboxw[8]), 
	.A(FE_PHN1256_prev_key1_reg_112_));
   XOR2X1 U1516 (.Y(n708), 
	.B(new_sboxw[14]), 
	.A(FE_PHN1313_prev_key1_reg_118_));
   XOR2X1 U1517 (.Y(n713), 
	.B(new_sboxw[9]), 
	.A(FE_PHN1236_prev_key1_reg_113_));
   XOR2X1 U1518 (.Y(n711), 
	.B(new_sboxw[11]), 
	.A(FE_PHN1244_prev_key1_reg_115_));
   XOR2X1 U1519 (.Y(n710), 
	.B(new_sboxw[12]), 
	.A(FE_PHN1249_prev_key1_reg_116_));
   XOR2X1 U1520 (.Y(n726), 
	.B(new_sboxw[28]), 
	.A(FE_PHN1225_prev_key1_reg_100_));
   XOR2X1 U1521 (.Y(n724), 
	.B(new_sboxw[30]), 
	.A(FE_PHN1220_prev_key1_reg_102_));
   XOR2X1 U1522 (.Y(n694), 
	.B(new_sboxw[22]), 
	.A(FE_PHN1989_rcon_reg_6_));
   AOI22X1 U1524 (.Y(n574), 
	.B1(n2652), 
	.B0(key[96]), 
	.A1(n730), 
	.A0(FE_OFN91_n690));
   AOI22X1 U1526 (.Y(n550), 
	.B1(n705), 
	.B0(FE_OFN91_n690), 
	.A1(n2640), 
	.A0(key[120]));
   XOR2X1 U1527 (.Y(n705), 
	.B(n706), 
	.A(FE_PHN1416_prev_key1_reg_120_));
   AOI22X1 U1529 (.Y(n544), 
	.B1(n693), 
	.B0(FE_OFN91_n690), 
	.A1(n2637), 
	.A0(key[126]));
   XOR2X1 U1530 (.Y(n693), 
	.B(n694), 
	.A(prev_key1_reg[126]));
   AOI22X1 U1532 (.Y(n545), 
	.B1(n695), 
	.B0(FE_OFN90_n690), 
	.A1(n2638), 
	.A0(key[125]));
   XOR2X1 U1533 (.Y(n695), 
	.B(n696), 
	.A(FE_PHN1391_prev_key1_reg_125_));
   AOI22X1 U1535 (.Y(n547), 
	.B1(n699), 
	.B0(FE_OFN90_n690), 
	.A1(n2639), 
	.A0(key[123]));
   XOR2X1 U1536 (.Y(n699), 
	.B(n700), 
	.A(FE_PHN1413_prev_key1_reg_123_));
   AOI22X1 U1538 (.Y(n549), 
	.B1(n703), 
	.B0(FE_OFN91_n690), 
	.A1(n2640), 
	.A0(key[121]));
   XOR2X1 U1539 (.Y(n703), 
	.B(n704), 
	.A(FE_PHN1395_prev_key1_reg_121_));
   XNOR2X1 U1540 (.Y(n806), 
	.B(n726), 
	.A(n866));
   XNOR2X1 U1541 (.Y(n866), 
	.B(FE_PHN1446_prev_key1_reg_68_), 
	.A(FE_PHN1053_prev_key1_reg_36_));
   XNOR2X1 U1542 (.Y(n805), 
	.B(n725), 
	.A(n864));
   XNOR2X1 U1543 (.Y(n864), 
	.B(FE_PHN1445_prev_key1_reg_69_), 
	.A(FE_PHN1056_prev_key1_reg_37_));
   XNOR2X1 U1544 (.Y(n804), 
	.B(n724), 
	.A(n862));
   XNOR2X1 U1545 (.Y(n862), 
	.B(prev_key1_reg[70]), 
	.A(FE_PHN1055_prev_key1_reg_38_));
   XNOR2X1 U1546 (.Y(n803), 
	.B(n723), 
	.A(n860));
   XNOR2X1 U1547 (.Y(n860), 
	.B(FE_PHN1406_prev_key1_reg_71_), 
	.A(FE_PHN1049_prev_key1_reg_39_));
   XNOR2X1 U1548 (.Y(n796), 
	.B(n716), 
	.A(n846));
   XNOR2X1 U1549 (.Y(n846), 
	.B(FE_PHN1402_prev_key1_reg_78_), 
	.A(prev_key1_reg[46]));
   XNOR2X1 U1550 (.Y(n794), 
	.B(n714), 
	.A(n842));
   XNOR2X1 U1551 (.Y(n842), 
	.B(FE_PHN1414_prev_key1_reg_80_), 
	.A(prev_key1_reg[48]));
   XNOR2X1 U1552 (.Y(n793), 
	.B(n713), 
	.A(n840));
   XNOR2X1 U1553 (.Y(n840), 
	.B(FE_PHN1425_prev_key1_reg_81_), 
	.A(FE_PHN1067_prev_key1_reg_49_));
   XNOR2X1 U1554 (.Y(n792), 
	.B(n712), 
	.A(n838));
   XNOR2X1 U1555 (.Y(n838), 
	.B(FE_PHN1405_prev_key1_reg_82_), 
	.A(FE_PHN1074_prev_key1_reg_50_));
   XNOR2X1 U1556 (.Y(n791), 
	.B(n711), 
	.A(n836));
   XNOR2X1 U1557 (.Y(n836), 
	.B(FE_PHN1388_prev_key1_reg_83_), 
	.A(FE_PHN1052_prev_key1_reg_51_));
   XNOR2X1 U1558 (.Y(n790), 
	.B(n710), 
	.A(n834));
   XNOR2X1 U1559 (.Y(n834), 
	.B(FE_PHN1375_prev_key1_reg_84_), 
	.A(FE_PHN1043_prev_key1_reg_52_));
   XNOR2X1 U1561 (.Y(n789), 
	.B(n709), 
	.A(n832));
   XNOR2X1 U1562 (.Y(n832), 
	.B(FE_PHN1412_prev_key1_reg_85_), 
	.A(FE_PHN1230_prev_key1_reg_53_));
   XNOR2X1 U1563 (.Y(n788), 
	.B(n708), 
	.A(n830));
   XNOR2X1 U1564 (.Y(n830), 
	.B(FE_PHN360_prev_key1_reg_86_), 
	.A(FE_PHN1050_prev_key1_reg_54_));
   XNOR2X1 U1565 (.Y(n787), 
	.B(n707), 
	.A(n828));
   XNOR2X1 U1566 (.Y(n828), 
	.B(FE_PHN359_prev_key1_reg_87_), 
	.A(FE_PHN1057_prev_key1_reg_55_));
   OAI2BB2X1 U1567 (.Y(n1254), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN571_n656), 
	.A1N(key_mem[1038]), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1568 (.Y(n1253), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN327_n655), 
	.A1N(FE_PHN1888_key_mem_1039_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1569 (.Y(n1251), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN570_n653), 
	.A1N(FE_PHN1840_key_mem_1041_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1570 (.Y(n1250), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN558_n652), 
	.A1N(FE_PHN1719_key_mem_1042_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1571 (.Y(n1249), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN569_n651), 
	.A1N(FE_PHN1833_key_mem_1043_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1572 (.Y(n1247), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN625_n649), 
	.A1N(FE_PHN1880_key_mem_1045_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1573 (.Y(n1246), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN564_n648), 
	.A1N(FE_PHN1905_key_mem_1046_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1574 (.Y(n1245), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN348_n647), 
	.A1N(FE_PHN1761_key_mem_1047_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1575 (.Y(n1126), 
	.B1(FE_OFN81_n672), 
	.B0(FE_PHN571_n656), 
	.A1N(FE_PHN798_key_mem_1166_), 
	.A0N(FE_OFN81_n672));
   OAI2BB2X1 U1576 (.Y(n1125), 
	.B1(FE_OFN81_n672), 
	.B0(FE_PHN327_n655), 
	.A1N(FE_PHN430_key_mem_1167_), 
	.A0N(FE_OFN81_n672));
   OAI2BB2X1 U1577 (.Y(n1123), 
	.B1(FE_OFN81_n672), 
	.B0(FE_PHN570_n653), 
	.A1N(FE_PHN1792_key_mem_1169_), 
	.A0N(FE_OFN81_n672));
   OAI2BB2X1 U1578 (.Y(n1122), 
	.B1(FE_OFN81_n672), 
	.B0(FE_PHN558_n652), 
	.A1N(FE_PHN582_key_mem_1170_), 
	.A0N(FE_OFN81_n672));
   OAI2BB2X1 U1579 (.Y(n1121), 
	.B1(FE_OFN81_n672), 
	.B0(FE_PHN569_n651), 
	.A1N(FE_PHN2839_key_mem_1171_), 
	.A0N(FE_OFN81_n672));
   OAI2BB2X1 U1580 (.Y(n1119), 
	.B1(FE_OFN81_n672), 
	.B0(FE_PHN625_n649), 
	.A1N(FE_PHN768_key_mem_1173_), 
	.A0N(FE_OFN81_n672));
   OAI2BB2X1 U1581 (.Y(n1118), 
	.B1(FE_OFN81_n672), 
	.B0(FE_PHN564_n648), 
	.A1N(FE_PHN1000_key_mem_1174_), 
	.A0N(FE_OFN81_n672));
   OAI2BB2X1 U1582 (.Y(n1117), 
	.B1(FE_OFN81_n672), 
	.B0(FE_PHN348_n647), 
	.A1N(FE_PHN585_key_mem_1175_), 
	.A0N(FE_OFN81_n672));
   OAI2BB2X1 U1583 (.Y(n1382), 
	.B1(FE_OFN76_n676), 
	.B0(FE_PHN571_n656), 
	.A1N(key_mem[910]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U1584 (.Y(n1381), 
	.B1(FE_OFN76_n676), 
	.B0(FE_PHN327_n655), 
	.A1N(key_mem[911]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U1585 (.Y(n1379), 
	.B1(FE_OFN76_n676), 
	.B0(FE_PHN570_n653), 
	.A1N(key_mem[913]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U1586 (.Y(n1378), 
	.B1(FE_OFN76_n676), 
	.B0(FE_PHN558_n652), 
	.A1N(key_mem[914]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U1587 (.Y(n1377), 
	.B1(FE_OFN76_n676), 
	.B0(FE_PHN569_n651), 
	.A1N(key_mem[915]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U1588 (.Y(n1375), 
	.B1(FE_OFN76_n676), 
	.B0(FE_PHN625_n649), 
	.A1N(key_mem[917]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U1589 (.Y(n1374), 
	.B1(FE_OFN76_n676), 
	.B0(FE_PHN564_n648), 
	.A1N(key_mem[918]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U1590 (.Y(n1373), 
	.B1(FE_OFN76_n676), 
	.B0(FE_PHN348_n647), 
	.A1N(key_mem[919]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U1591 (.Y(n998), 
	.B1(FE_OFN85_n1), 
	.B0(FE_PHN571_n656), 
	.A1N(key_mem[1294]), 
	.A0N(FE_OFN85_n1));
   OAI2BB2X1 U1592 (.Y(n997), 
	.B1(FE_OFN85_n1), 
	.B0(FE_PHN327_n655), 
	.A1N(FE_PHN2840_key_mem_1295_), 
	.A0N(FE_OFN85_n1));
   OAI2BB2X1 U1593 (.Y(n995), 
	.B1(FE_OFN85_n1), 
	.B0(FE_PHN570_n653), 
	.A1N(FE_PHN2837_key_mem_1297_), 
	.A0N(FE_OFN85_n1));
   OAI2BB2X1 U1594 (.Y(n994), 
	.B1(n1), 
	.B0(FE_PHN558_n652), 
	.A1N(FE_PHN2823_key_mem_1298_), 
	.A0N(n1));
   OAI2BB2X1 U1595 (.Y(n993), 
	.B1(FE_OFN85_n1), 
	.B0(FE_PHN569_n651), 
	.A1N(FE_PHN3435_key_mem_1299_), 
	.A0N(FE_OFN85_n1));
   OAI2BB2X1 U1596 (.Y(n991), 
	.B1(FE_OFN85_n1), 
	.B0(FE_PHN625_n649), 
	.A1N(key_mem[1301]), 
	.A0N(FE_OFN85_n1));
   OAI2BB2X1 U1597 (.Y(n990), 
	.B1(FE_OFN85_n1), 
	.B0(FE_PHN564_n648), 
	.A1N(FE_PHN2835_key_mem_1302_), 
	.A0N(FE_OFN85_n1));
   OAI2BB2X1 U1598 (.Y(n989), 
	.B1(FE_OFN85_n1), 
	.B0(FE_PHN348_n647), 
	.A1N(FE_PHN3094_key_mem_1303_), 
	.A0N(FE_OFN85_n1));
   OAI2BB2X1 U1599 (.Y(n1365), 
	.B1(FE_OFN76_n676), 
	.B0(FE_PHN401_n639), 
	.A1N(key_mem[927]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U1600 (.Y(n1237), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN401_n639), 
	.A1N(FE_PHN1864_key_mem_1055_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1601 (.Y(n1109), 
	.B1(FE_OFN81_n672), 
	.B0(FE_PHN401_n639), 
	.A1N(FE_PHN3319_key_mem_1183_), 
	.A0N(FE_OFN81_n672));
   OAI2BB2X1 U1602 (.Y(n981), 
	.B1(FE_OFN85_n1), 
	.B0(FE_PHN401_n639), 
	.A1N(FE_PHN1834_key_mem_1311_), 
	.A0N(FE_OFN85_n1));
   OAI2BB2X1 U1603 (.Y(n1333), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN423_n607), 
	.A1N(key_mem[959]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1604 (.Y(n1205), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN423_n607), 
	.A1N(key_mem[1087]), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U1605 (.Y(n1077), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN423_n607), 
	.A1N(FE_PHN1700_key_mem_1215_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1606 (.Y(n949), 
	.B1(FE_OFN88_n1), 
	.B0(FE_PHN423_n607), 
	.A1N(key_mem[1343]), 
	.A0N(FE_OFN88_n1));
   OAI2BB2X1 U1607 (.Y(n1301), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN342_n575), 
	.A1N(key_mem[991]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1608 (.Y(n1173), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN342_n575), 
	.A1N(FE_PHN1817_key_mem_1119_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1609 (.Y(n1045), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN342_n575), 
	.A1N(FE_PHN811_key_mem_1247_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1610 (.Y(n917), 
	.B1(n2623), 
	.B0(FE_PHN342_n575), 
	.A1N(FE_PHN2833_key_mem_1375_), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U1611 (.Y(n1269), 
	.B1(FE_OFN76_n676), 
	.B0(FE_PHN622_n543), 
	.A1N(key_mem[1023]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U1612 (.Y(n1141), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN622_n543), 
	.A1N(FE_PHN1884_key_mem_1151_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1613 (.Y(n1013), 
	.B1(FE_OFN81_n672), 
	.B0(FE_PHN622_n543), 
	.A1N(FE_PHN3091_key_mem_1279_), 
	.A0N(FE_OFN81_n672));
   OAI2BB2X1 U1614 (.Y(n885), 
	.B1(n1), 
	.B0(FE_PHN622_n543), 
	.A1N(FE_PHN3444_key_mem_1407_), 
	.A0N(FE_OFN85_n1));
   OAI2BB2X1 U1615 (.Y(n1372), 
	.B1(FE_OFN76_n676), 
	.B0(FE_PHN406_n646), 
	.A1N(key_mem[920]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U1616 (.Y(n1244), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN406_n646), 
	.A1N(key_mem[1048]), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1617 (.Y(n1116), 
	.B1(FE_OFN81_n672), 
	.B0(FE_PHN406_n646), 
	.A1N(FE_PHN819_key_mem_1176_), 
	.A0N(FE_OFN81_n672));
   OAI2BB2X1 U1618 (.Y(n988), 
	.B1(FE_OFN85_n1), 
	.B0(FE_PHN406_n646), 
	.A1N(FE_PHN2827_key_mem_1304_), 
	.A0N(FE_OFN85_n1));
   OAI2BB2X1 U1619 (.Y(n1340), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN404_n614), 
	.A1N(key_mem[952]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1620 (.Y(n1212), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN404_n614), 
	.A1N(FE_PHN1730_key_mem_1080_), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1621 (.Y(n1084), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN404_n614), 
	.A1N(FE_PHN786_key_mem_1208_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1622 (.Y(n956), 
	.B1(FE_OFN87_n1), 
	.B0(FE_PHN404_n614), 
	.A1N(key_mem[1336]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U1623 (.Y(n1308), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN347_n582), 
	.A1N(key_mem[984]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1624 (.Y(n1180), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN347_n582), 
	.A1N(FE_PHN1860_key_mem_1112_), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U1625 (.Y(n1052), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN347_n582), 
	.A1N(FE_PHN817_key_mem_1240_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1626 (.Y(n924), 
	.B1(n2624), 
	.B0(FE_PHN347_n582), 
	.A1N(FE_PHN2830_key_mem_1368_), 
	.A0N(n1));
   OAI2BB2X1 U1627 (.Y(n1276), 
	.B1(FE_OFN76_n676), 
	.B0(FE_PHN568_n550), 
	.A1N(key_mem[1016]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U1628 (.Y(n1148), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN568_n550), 
	.A1N(FE_PHN1858_key_mem_1144_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1629 (.Y(n1020), 
	.B1(n672), 
	.B0(FE_PHN568_n550), 
	.A1N(FE_PHN1899_key_mem_1272_), 
	.A0N(n672));
   OAI2BB2X1 U1630 (.Y(n892), 
	.B1(FE_OFN85_n1), 
	.B0(FE_PHN568_n550), 
	.A1N(FE_PHN3229_key_mem_1400_), 
	.A0N(FE_OFN85_n1));
   OAI2BB2X1 U1631 (.Y(n1366), 
	.B1(FE_OFN76_n676), 
	.B0(FE_PHN408_n640), 
	.A1N(key_mem[926]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U1632 (.Y(n1238), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN408_n640), 
	.A1N(FE_PHN1769_key_mem_1054_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1633 (.Y(n1110), 
	.B1(FE_OFN81_n672), 
	.B0(FE_PHN408_n640), 
	.A1N(FE_PHN808_key_mem_1182_), 
	.A0N(FE_OFN81_n672));
   OAI2BB2X1 U1634 (.Y(n982), 
	.B1(FE_OFN85_n1), 
	.B0(FE_PHN408_n640), 
	.A1N(key_mem[1310]), 
	.A0N(FE_OFN85_n1));
   OAI2BB2X1 U1635 (.Y(n1334), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN422_n608), 
	.A1N(key_mem[958]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1636 (.Y(n1206), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN422_n608), 
	.A1N(key_mem[1086]), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1637 (.Y(n1078), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN422_n608), 
	.A1N(FE_PHN800_key_mem_1214_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1638 (.Y(n950), 
	.B1(FE_OFN88_n1), 
	.B0(FE_PHN422_n608), 
	.A1N(key_mem[1342]), 
	.A0N(FE_OFN88_n1));
   OAI2BB2X1 U1639 (.Y(n1302), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN344_n576), 
	.A1N(key_mem[990]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1640 (.Y(n1174), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN344_n576), 
	.A1N(FE_PHN1803_key_mem_1118_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1641 (.Y(n1046), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN344_n576), 
	.A1N(FE_PHN794_key_mem_1246_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1642 (.Y(n918), 
	.B1(n2623), 
	.B0(FE_PHN344_n576), 
	.A1N(key_mem[1374]), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U1643 (.Y(n1270), 
	.B1(FE_OFN76_n676), 
	.B0(FE_PHN623_n544), 
	.A1N(key_mem[1022]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U1644 (.Y(n1142), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN623_n544), 
	.A1N(FE_PHN1814_key_mem_1150_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1645 (.Y(n1014), 
	.B1(FE_OFN81_n672), 
	.B0(FE_PHN623_n544), 
	.A1N(FE_PHN1766_key_mem_1278_), 
	.A0N(FE_OFN81_n672));
   OAI2BB2X1 U1646 (.Y(n886), 
	.B1(FE_OFN85_n1), 
	.B0(FE_PHN623_n544), 
	.A1N(key_mem[1406]), 
	.A0N(FE_OFN85_n1));
   OAI2BB2X1 U1647 (.Y(n1367), 
	.B1(n676), 
	.B0(FE_PHN400_n641), 
	.A1N(key_mem[925]), 
	.A0N(n676));
   OAI2BB2X1 U1648 (.Y(n1239), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN400_n641), 
	.A1N(FE_PHN1868_key_mem_1053_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1649 (.Y(n1111), 
	.B1(n672), 
	.B0(FE_PHN400_n641), 
	.A1N(key_mem[1181]), 
	.A0N(n672));
   OAI2BB2X1 U1650 (.Y(n983), 
	.B1(FE_OFN87_n1), 
	.B0(FE_PHN400_n641), 
	.A1N(key_mem[1309]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U1651 (.Y(n1335), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN393_n609), 
	.A1N(key_mem[957]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1652 (.Y(n1207), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN393_n609), 
	.A1N(FE_PHN1856_key_mem_1085_), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1653 (.Y(n1079), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN393_n609), 
	.A1N(FE_PHN782_key_mem_1213_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1654 (.Y(n951), 
	.B1(FE_OFN89_n1), 
	.B0(FE_PHN393_n609), 
	.A1N(key_mem[1341]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U1655 (.Y(n1303), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN343_n577), 
	.A1N(key_mem[989]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1656 (.Y(n1175), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN343_n577), 
	.A1N(key_mem[1117]), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U1657 (.Y(n1047), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN343_n577), 
	.A1N(FE_PHN773_key_mem_1245_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1658 (.Y(n919), 
	.B1(n2623), 
	.B0(FE_PHN343_n577), 
	.A1N(key_mem[1373]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U1659 (.Y(n1271), 
	.B1(n676), 
	.B0(FE_PHN551_n545), 
	.A1N(key_mem[1021]), 
	.A0N(n676));
   OAI2BB2X1 U1660 (.Y(n1143), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN551_n545), 
	.A1N(key_mem[1149]), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1661 (.Y(n1015), 
	.B1(n672), 
	.B0(FE_PHN551_n545), 
	.A1N(FE_PHN792_key_mem_1277_), 
	.A0N(n672));
   OAI2BB2X1 U1662 (.Y(n887), 
	.B1(FE_OFN87_n1), 
	.B0(FE_PHN551_n545), 
	.A1N(key_mem[1405]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U1663 (.Y(n1368), 
	.B1(n676), 
	.B0(FE_PHN397_n642), 
	.A1N(key_mem[924]), 
	.A0N(n676));
   OAI2BB2X1 U1664 (.Y(n1240), 
	.B1(n674), 
	.B0(FE_PHN397_n642), 
	.A1N(key_mem[1052]), 
	.A0N(n674));
   OAI2BB2X1 U1665 (.Y(n1112), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN397_n642), 
	.A1N(key_mem[1180]), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1666 (.Y(n984), 
	.B1(FE_OFN87_n1), 
	.B0(FE_PHN397_n642), 
	.A1N(key_mem[1308]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U1667 (.Y(n1336), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN392_n610), 
	.A1N(key_mem[956]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1668 (.Y(n1208), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN392_n610), 
	.A1N(FE_PHN1835_key_mem_1084_), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1669 (.Y(n1080), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN392_n610), 
	.A1N(FE_PHN797_key_mem_1212_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1670 (.Y(n952), 
	.B1(FE_OFN89_n1), 
	.B0(FE_PHN392_n610), 
	.A1N(key_mem[1340]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U1671 (.Y(n1304), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN345_n578), 
	.A1N(key_mem[988]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1672 (.Y(n1176), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN345_n578), 
	.A1N(FE_PHN1843_key_mem_1116_), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1673 (.Y(n1048), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN345_n578), 
	.A1N(key_mem[1244]), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1674 (.Y(n920), 
	.B1(n2623), 
	.B0(FE_PHN345_n578), 
	.A1N(FE_PHN788_key_mem_1372_), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U1675 (.Y(n1272), 
	.B1(n676), 
	.B0(FE_PHN548_n546), 
	.A1N(key_mem[1020]), 
	.A0N(n676));
   OAI2BB2X1 U1676 (.Y(n1144), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN548_n546), 
	.A1N(FE_PHN1808_key_mem_1148_), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U1677 (.Y(n1016), 
	.B1(n672), 
	.B0(FE_PHN548_n546), 
	.A1N(FE_PHN780_key_mem_1276_), 
	.A0N(n672));
   OAI2BB2X1 U1678 (.Y(n888), 
	.B1(FE_OFN87_n1), 
	.B0(FE_PHN548_n546), 
	.A1N(key_mem[1404]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U1679 (.Y(n1369), 
	.B1(n676), 
	.B0(FE_PHN399_n643), 
	.A1N(key_mem[923]), 
	.A0N(n676));
   OAI2BB2X1 U1680 (.Y(n1241), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN399_n643), 
	.A1N(FE_PHN1784_key_mem_1051_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1681 (.Y(n1113), 
	.B1(n672), 
	.B0(FE_PHN399_n643), 
	.A1N(FE_PHN760_key_mem_1179_), 
	.A0N(n672));
   OAI2BB2X1 U1682 (.Y(n985), 
	.B1(n1), 
	.B0(FE_PHN399_n643), 
	.A1N(key_mem[1307]), 
	.A0N(n1));
   OAI2BB2X1 U1683 (.Y(n1337), 
	.B1(n676), 
	.B0(FE_PHN386_n611), 
	.A1N(key_mem[955]), 
	.A0N(n676));
   OAI2BB2X1 U1684 (.Y(n1209), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN386_n611), 
	.A1N(FE_PHN1857_key_mem_1083_), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U1685 (.Y(n1081), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN386_n611), 
	.A1N(FE_PHN765_key_mem_1211_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1686 (.Y(n953), 
	.B1(FE_OFN87_n1), 
	.B0(FE_PHN386_n611), 
	.A1N(key_mem[1339]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U1687 (.Y(n1305), 
	.B1(n676), 
	.B0(FE_PHN346_n579), 
	.A1N(key_mem[987]), 
	.A0N(n676));
   OAI2BB2X1 U1688 (.Y(n1177), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN346_n579), 
	.A1N(FE_PHN1823_key_mem_1115_), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U1689 (.Y(n1049), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN346_n579), 
	.A1N(FE_PHN771_key_mem_1243_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1691 (.Y(n921), 
	.B1(n2623), 
	.B0(FE_PHN346_n579), 
	.A1N(key_mem[1371]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U1692 (.Y(n1273), 
	.B1(n676), 
	.B0(FE_PHN544_n547), 
	.A1N(key_mem[1019]), 
	.A0N(n676));
   OAI2BB2X1 U1693 (.Y(n1145), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN544_n547), 
	.A1N(FE_PHN1805_key_mem_1147_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1694 (.Y(n1017), 
	.B1(n672), 
	.B0(FE_PHN544_n547), 
	.A1N(key_mem[1275]), 
	.A0N(n672));
   OAI2BB2X1 U1695 (.Y(n889), 
	.B1(FE_OFN87_n1), 
	.B0(FE_PHN544_n547), 
	.A1N(key_mem[1403]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U1696 (.Y(n1338), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN326_n612), 
	.A1N(key_mem[954]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1697 (.Y(n1210), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN326_n612), 
	.A1N(FE_PHN1930_key_mem_1082_), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U1698 (.Y(n1082), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN326_n612), 
	.A1N(key_mem[1210]), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1699 (.Y(n954), 
	.B1(FE_OFN87_n1), 
	.B0(FE_PHN326_n612), 
	.A1N(key_mem[1338]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U1700 (.Y(n1306), 
	.B1(n676), 
	.B0(FE_PHN547_n580), 
	.A1N(key_mem[986]), 
	.A0N(n676));
   OAI2BB2X1 U1701 (.Y(n1178), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN547_n580), 
	.A1N(FE_PHN1885_key_mem_1114_), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U1702 (.Y(n1050), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN547_n580), 
	.A1N(FE_PHN767_key_mem_1242_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1703 (.Y(n922), 
	.B1(n2624), 
	.B0(FE_PHN547_n580), 
	.A1N(key_mem[1370]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U1704 (.Y(n1274), 
	.B1(n676), 
	.B0(FE_PHN418_n548), 
	.A1N(key_mem[1018]), 
	.A0N(n676));
   OAI2BB2X1 U1705 (.Y(n1146), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN418_n548), 
	.A1N(key_mem[1146]), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1706 (.Y(n1018), 
	.B1(n672), 
	.B0(FE_PHN418_n548), 
	.A1N(FE_PHN766_key_mem_1274_), 
	.A0N(n672));
   OAI2BB2X1 U1707 (.Y(n890), 
	.B1(FE_OFN87_n1), 
	.B0(FE_PHN418_n548), 
	.A1N(key_mem[1402]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U1708 (.Y(n1371), 
	.B1(FE_OFN76_n676), 
	.B0(FE_PHN407_n645), 
	.A1N(key_mem[921]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U1709 (.Y(n1243), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN407_n645), 
	.A1N(FE_PHN1876_key_mem_1049_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1710 (.Y(n1115), 
	.B1(n672), 
	.B0(FE_PHN407_n645), 
	.A1N(FE_PHN791_key_mem_1177_), 
	.A0N(n672));
   OAI2BB2X1 U1711 (.Y(n987), 
	.B1(n1), 
	.B0(FE_PHN407_n645), 
	.A1N(FE_PHN2829_key_mem_1305_), 
	.A0N(n1));
   OAI2BB2X1 U1712 (.Y(n1339), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN405_n613), 
	.A1N(key_mem[953]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1713 (.Y(n1211), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN405_n613), 
	.A1N(FE_PHN1783_key_mem_1081_), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1714 (.Y(n1083), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN405_n613), 
	.A1N(FE_PHN783_key_mem_1209_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1715 (.Y(n955), 
	.B1(FE_OFN89_n1), 
	.B0(FE_PHN405_n613), 
	.A1N(key_mem[1337]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U1716 (.Y(n1307), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN349_n581), 
	.A1N(key_mem[985]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1717 (.Y(n1179), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN349_n581), 
	.A1N(FE_PHN1818_key_mem_1113_), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1718 (.Y(n1051), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN349_n581), 
	.A1N(FE_PHN770_key_mem_1241_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1719 (.Y(n923), 
	.B1(n2624), 
	.B0(FE_PHN349_n581), 
	.A1N(key_mem[1369]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U1720 (.Y(n1275), 
	.B1(FE_OFN76_n676), 
	.B0(FE_PHN567_n549), 
	.A1N(key_mem[1017]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U1721 (.Y(n1147), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN567_n549), 
	.A1N(FE_PHN1762_key_mem_1145_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1722 (.Y(n1019), 
	.B1(n672), 
	.B0(FE_PHN567_n549), 
	.A1N(FE_PHN802_key_mem_1273_), 
	.A0N(n672));
   OAI2BB2X1 U1723 (.Y(n891), 
	.B1(n1), 
	.B0(FE_PHN567_n549), 
	.A1N(FE_PHN2834_key_mem_1401_), 
	.A0N(n1));
   OAI2BB2X1 U1724 (.Y(n1268), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN553_n670), 
	.A1N(key_mem[1024]), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1725 (.Y(n1267), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN537_n669), 
	.A1N(FE_PHN1882_key_mem_1025_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1726 (.Y(n1266), 
	.B1(n674), 
	.B0(FE_PHN550_n668), 
	.A1N(FE_PHN3239_key_mem_1026_), 
	.A0N(n674));
   OAI2BB2X1 U1727 (.Y(n1265), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN563_n667), 
	.A1N(key_mem[1027]), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1728 (.Y(n1264), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN562_n666), 
	.A1N(FE_PHN1853_key_mem_1028_), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U1729 (.Y(n1263), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN566_n665), 
	.A1N(FE_PHN1892_key_mem_1029_), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U1730 (.Y(n1262), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN572_n664), 
	.A1N(FE_PHN1862_key_mem_1030_), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U1731 (.Y(n1261), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN324_n663), 
	.A1N(FE_PHN1760_key_mem_1031_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1732 (.Y(n1260), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN325_n662), 
	.A1N(FE_PHN1713_key_mem_1032_), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U1733 (.Y(n1259), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN323_n661), 
	.A1N(FE_PHN2838_key_mem_1033_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1734 (.Y(n1258), 
	.B1(n674), 
	.B0(FE_PHN541_n660), 
	.A1N(FE_PHN3303_key_mem_1034_), 
	.A0N(n674));
   OAI2BB2X1 U1735 (.Y(n1257), 
	.B1(n674), 
	.B0(FE_PHN554_n659), 
	.A1N(key_mem[1035]), 
	.A0N(n674));
   OAI2BB2X1 U1736 (.Y(n1256), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN560_n658), 
	.A1N(FE_PHN1811_key_mem_1036_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1737 (.Y(n1255), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN552_n657), 
	.A1N(FE_PHN1788_key_mem_1037_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1738 (.Y(n1252), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN573_n654), 
	.A1N(FE_PHN1881_key_mem_1040_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1739 (.Y(n1248), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN579_n650), 
	.A1N(FE_PHN1894_key_mem_1044_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1740 (.Y(n1236), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN383_n638), 
	.A1N(key_mem[1056]), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1741 (.Y(n1235), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN380_n637), 
	.A1N(FE_PHN1832_key_mem_1057_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1742 (.Y(n1234), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN381_n636), 
	.A1N(FE_PHN1743_key_mem_1058_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1743 (.Y(n1233), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN379_n635), 
	.A1N(FE_PHN1839_key_mem_1059_), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U1744 (.Y(n1232), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN394_n634), 
	.A1N(FE_PHN1872_key_mem_1060_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1745 (.Y(n1231), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN391_n633), 
	.A1N(FE_PHN1873_key_mem_1061_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1746 (.Y(n1230), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN396_n632), 
	.A1N(key_mem[1062]), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1747 (.Y(n1229), 
	.B1(FE_OFN96_n674), 
	.B0(n631), 
	.A1N(FE_PHN954_key_mem_1063_), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1748 (.Y(n1228), 
	.B1(FE_OFN96_n674), 
	.B0(n630), 
	.A1N(FE_PHN1852_key_mem_1064_), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1749 (.Y(n1227), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN705_n629), 
	.A1N(key_mem[1065]), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1750 (.Y(n1226), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN390_n628), 
	.A1N(FE_PHN1813_key_mem_1066_), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1751 (.Y(n1225), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN398_n627), 
	.A1N(key_mem[1067]), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1752 (.Y(n1224), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN388_n626), 
	.A1N(FE_PHN1891_key_mem_1068_), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1753 (.Y(n1223), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN387_n625), 
	.A1N(FE_PHN1867_key_mem_1069_), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1754 (.Y(n1222), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN409_n624), 
	.A1N(FE_PHN1758_key_mem_1070_), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1755 (.Y(n1221), 
	.B1(FE_OFN96_n674), 
	.B0(n623), 
	.A1N(FE_PHN1889_key_mem_1071_), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1756 (.Y(n1220), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN403_n622), 
	.A1N(FE_PHN1861_key_mem_1072_), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1757 (.Y(n1219), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN402_n621), 
	.A1N(key_mem[1073]), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1758 (.Y(n1218), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN384_n620), 
	.A1N(FE_PHN1773_key_mem_1074_), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1759 (.Y(n1217), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN382_n619), 
	.A1N(FE_PHN1712_key_mem_1075_), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U1760 (.Y(n1215), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN385_n617), 
	.A1N(FE_PHN1789_key_mem_1077_), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1761 (.Y(n1214), 
	.B1(FE_OFN96_n674), 
	.B0(n616), 
	.A1N(FE_PHN1866_key_mem_1078_), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1762 (.Y(n1213), 
	.B1(FE_OFN96_n674), 
	.B0(n615), 
	.A1N(FE_PHN1829_key_mem_1079_), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1763 (.Y(n1204), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN540_n606), 
	.A1N(FE_PHN1869_key_mem_1088_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1764 (.Y(n1203), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN555_n605), 
	.A1N(FE_PHN1701_key_mem_1089_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1765 (.Y(n1202), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN538_n604), 
	.A1N(FE_PHN1830_key_mem_1090_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1766 (.Y(n1201), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN546_n603), 
	.A1N(key_mem[1091]), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1767 (.Y(n1200), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN557_n602), 
	.A1N(FE_PHN1841_key_mem_1092_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1768 (.Y(n1199), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN561_n601), 
	.A1N(FE_PHN1790_key_mem_1093_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1769 (.Y(n1197), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN545_n599), 
	.A1N(FE_PHN1778_key_mem_1095_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1770 (.Y(n1196), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN559_n598), 
	.A1N(key_mem[1096]), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1771 (.Y(n1195), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN416_n597), 
	.A1N(FE_PHN1799_key_mem_1097_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1772 (.Y(n1194), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN565_n596), 
	.A1N(FE_PHN1756_key_mem_1098_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1773 (.Y(n1193), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN556_n595), 
	.A1N(FE_PHN1859_key_mem_1099_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1774 (.Y(n1192), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN575_n594), 
	.A1N(FE_PHN1887_key_mem_1100_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1775 (.Y(n1191), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN577_n593), 
	.A1N(FE_PHN1893_key_mem_1101_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1776 (.Y(n1190), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN420_n592), 
	.A1N(key_mem[1102]), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1777 (.Y(n1189), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN417_n591), 
	.A1N(FE_PHN1855_key_mem_1103_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1778 (.Y(n1186), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN543_n588), 
	.A1N(FE_PHN1871_key_mem_1106_), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U1779 (.Y(n1185), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN549_n587), 
	.A1N(key_mem[1107]), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U1780 (.Y(n1183), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN539_n585), 
	.A1N(FE_PHN1787_key_mem_1109_), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1781 (.Y(n1182), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN576_n584), 
	.A1N(key_mem[1110]), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U1782 (.Y(n1181), 
	.B1(n674), 
	.B0(FE_PHN574_n583), 
	.A1N(key_mem[1111]), 
	.A0N(n674));
   OAI2BB2X1 U1783 (.Y(n1172), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN609_n574), 
	.A1N(FE_PHN1740_key_mem_1120_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1784 (.Y(n1169), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN606_n571), 
	.A1N(FE_PHN1781_key_mem_1123_), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U1785 (.Y(n1164), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN607_n566), 
	.A1N(FE_PHN1816_key_mem_1128_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U1786 (.Y(n1163), 
	.B1(FE_OFN94_n674), 
	.B0(n565), 
	.A1N(key_mem[1129]), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1787 (.Y(n1162), 
	.B1(n674), 
	.B0(FE_PHN608_n564), 
	.A1N(FE_PHN3307_key_mem_1130_), 
	.A0N(n674));
   OAI2BB2X1 U1788 (.Y(n1161), 
	.B1(n674), 
	.B0(FE_PHN615_n563), 
	.A1N(key_mem[1131]), 
	.A0N(n674));
   OAI2BB2X1 U1789 (.Y(n1159), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN621_n561), 
	.A1N(FE_PHN1822_key_mem_1133_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1790 (.Y(n1157), 
	.B1(FE_OFN94_n674), 
	.B0(n559), 
	.A1N(FE_PHN1791_key_mem_1135_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U1791 (.Y(n1140), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN553_n670), 
	.A1N(FE_PHN1734_key_mem_1152_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1792 (.Y(n1139), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN537_n669), 
	.A1N(FE_PHN1883_key_mem_1153_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1793 (.Y(n1138), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN550_n668), 
	.A1N(FE_PHN357_key_mem_1154_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1794 (.Y(n1137), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN563_n667), 
	.A1N(FE_PHN1023_key_mem_1155_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1795 (.Y(n1136), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN562_n666), 
	.A1N(FE_PHN775_key_mem_1156_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1796 (.Y(n1135), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN566_n665), 
	.A1N(FE_PHN989_key_mem_1157_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1797 (.Y(n1134), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN572_n664), 
	.A1N(FE_PHN980_key_mem_1158_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1798 (.Y(n1133), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN324_n663), 
	.A1N(FE_PHN584_key_mem_1159_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1799 (.Y(n1132), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN325_n662), 
	.A1N(key_mem[1160]), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1800 (.Y(n1131), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN323_n661), 
	.A1N(FE_PHN587_key_mem_1161_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1801 (.Y(n1130), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN541_n660), 
	.A1N(FE_PHN429_key_mem_1162_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1802 (.Y(n1129), 
	.B1(n672), 
	.B0(FE_PHN554_n659), 
	.A1N(FE_PHN974_key_mem_1163_), 
	.A0N(n672));
   OAI2BB2X1 U1803 (.Y(n1128), 
	.B1(n672), 
	.B0(FE_PHN560_n658), 
	.A1N(key_mem[1164]), 
	.A0N(n672));
   OAI2BB2X1 U1804 (.Y(n1127), 
	.B1(n672), 
	.B0(FE_PHN552_n657), 
	.A1N(key_mem[1165]), 
	.A0N(n672));
   OAI2BB2X1 U1805 (.Y(n1124), 
	.B1(FE_OFN81_n672), 
	.B0(FE_PHN573_n654), 
	.A1N(key_mem[1168]), 
	.A0N(FE_OFN81_n672));
   OAI2BB2X1 U1806 (.Y(n1120), 
	.B1(FE_OFN81_n672), 
	.B0(FE_PHN579_n650), 
	.A1N(FE_PHN698_key_mem_1172_), 
	.A0N(FE_OFN81_n672));
   OAI2BB2X1 U1807 (.Y(n1108), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN383_n638), 
	.A1N(FE_PHN426_key_mem_1184_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1808 (.Y(n1107), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN380_n637), 
	.A1N(key_mem[1185]), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1809 (.Y(n1106), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN381_n636), 
	.A1N(FE_PHN1015_key_mem_1186_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1810 (.Y(n1105), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN379_n635), 
	.A1N(key_mem[1187]), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1811 (.Y(n1104), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN394_n634), 
	.A1N(FE_PHN1720_key_mem_1188_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1812 (.Y(n1103), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN391_n633), 
	.A1N(FE_PHN1083_key_mem_1189_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1813 (.Y(n1102), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN396_n632), 
	.A1N(key_mem[1190]), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1814 (.Y(n1101), 
	.B1(FE_OFN82_n672), 
	.B0(n631), 
	.A1N(FE_PHN1800_key_mem_1191_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1815 (.Y(n1100), 
	.B1(FE_OFN82_n672), 
	.B0(n630), 
	.A1N(FE_PHN1005_key_mem_1192_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1816 (.Y(n1099), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN705_n629), 
	.A1N(FE_PHN1029_key_mem_1193_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1817 (.Y(n1098), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN390_n628), 
	.A1N(FE_PHN696_key_mem_1194_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1818 (.Y(n1097), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN398_n627), 
	.A1N(FE_PHN943_key_mem_1195_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1820 (.Y(n1096), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN388_n626), 
	.A1N(FE_PHN929_key_mem_1196_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1821 (.Y(n1095), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN387_n625), 
	.A1N(key_mem[1197]), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1822 (.Y(n1094), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN409_n624), 
	.A1N(FE_PHN955_key_mem_1198_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1823 (.Y(n1093), 
	.B1(FE_OFN82_n672), 
	.B0(n623), 
	.A1N(FE_PHN1008_key_mem_1199_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1824 (.Y(n1092), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN403_n622), 
	.A1N(FE_PHN953_key_mem_1200_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1825 (.Y(n1091), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN402_n621), 
	.A1N(FE_PHN958_key_mem_1201_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1826 (.Y(n1090), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN384_n620), 
	.A1N(FE_PHN992_key_mem_1202_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1827 (.Y(n1089), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN382_n619), 
	.A1N(FE_PHN942_key_mem_1203_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1828 (.Y(n1087), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN385_n617), 
	.A1N(FE_PHN1024_key_mem_1205_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1829 (.Y(n1086), 
	.B1(FE_OFN80_n672), 
	.B0(n616), 
	.A1N(FE_PHN1021_key_mem_1206_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1830 (.Y(n1085), 
	.B1(FE_OFN80_n672), 
	.B0(n615), 
	.A1N(FE_PHN1917_key_mem_1207_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1831 (.Y(n1076), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN540_n606), 
	.A1N(key_mem[1216]), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1832 (.Y(n1075), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN555_n605), 
	.A1N(key_mem[1217]), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1833 (.Y(n1074), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN538_n604), 
	.A1N(FE_PHN785_key_mem_1218_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1834 (.Y(n1073), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN546_n603), 
	.A1N(FE_PHN1006_key_mem_1219_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1835 (.Y(n1072), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN557_n602), 
	.A1N(FE_PHN977_key_mem_1220_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1836 (.Y(n1071), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN561_n601), 
	.A1N(key_mem[1221]), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1837 (.Y(n1069), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN545_n599), 
	.A1N(FE_PHN689_key_mem_1223_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1838 (.Y(n1068), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN559_n598), 
	.A1N(FE_PHN431_key_mem_1224_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1839 (.Y(n1067), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN416_n597), 
	.A1N(FE_PHN594_key_mem_1225_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1840 (.Y(n1066), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN565_n596), 
	.A1N(FE_PHN692_key_mem_1226_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1841 (.Y(n1065), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN556_n595), 
	.A1N(FE_PHN975_key_mem_1227_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1842 (.Y(n1064), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN575_n594), 
	.A1N(FE_PHN960_key_mem_1228_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1843 (.Y(n1063), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN577_n593), 
	.A1N(FE_PHN934_key_mem_1229_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1844 (.Y(n1062), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN420_n592), 
	.A1N(FE_PHN591_key_mem_1230_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1845 (.Y(n1061), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN417_n591), 
	.A1N(FE_PHN949_key_mem_1231_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1846 (.Y(n1058), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN543_n588), 
	.A1N(FE_PHN777_key_mem_1234_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1847 (.Y(n1057), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN549_n587), 
	.A1N(FE_PHN972_key_mem_1235_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1848 (.Y(n1055), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN539_n585), 
	.A1N(key_mem[1237]), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1849 (.Y(n1054), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN576_n584), 
	.A1N(FE_PHN936_key_mem_1238_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1850 (.Y(n1053), 
	.B1(n672), 
	.B0(FE_PHN574_n583), 
	.A1N(FE_PHN776_key_mem_1239_), 
	.A0N(n672));
   OAI2BB2X1 U1851 (.Y(n1044), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN609_n574), 
	.A1N(FE_PHN691_key_mem_1248_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1852 (.Y(n1041), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN606_n571), 
	.A1N(key_mem[1251]), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U1853 (.Y(n1036), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN607_n566), 
	.A1N(FE_PHN432_key_mem_1256_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U1854 (.Y(n1035), 
	.B1(n672), 
	.B0(n565), 
	.A1N(FE_PHN583_key_mem_1257_), 
	.A0N(n672));
   OAI2BB2X1 U1855 (.Y(n1034), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN608_n564), 
	.A1N(FE_PHN427_key_mem_1258_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1856 (.Y(n1033), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN615_n563), 
	.A1N(FE_PHN1009_key_mem_1259_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U1857 (.Y(n1031), 
	.B1(n672), 
	.B0(FE_PHN621_n561), 
	.A1N(FE_PHN981_key_mem_1261_), 
	.A0N(n672));
   OAI2BB2X1 U1858 (.Y(n1029), 
	.B1(FE_OFN81_n672), 
	.B0(n559), 
	.A1N(FE_PHN2842_key_mem_1263_), 
	.A0N(FE_OFN81_n672));
   OAI2BB2X1 U1859 (.Y(n1396), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN553_n670), 
	.A1N(key_mem[896]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1860 (.Y(n1395), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN537_n669), 
	.A1N(key_mem[897]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1861 (.Y(n1394), 
	.B1(n676), 
	.B0(FE_PHN550_n668), 
	.A1N(FE_PHN3434_key_mem_898_), 
	.A0N(n676));
   OAI2BB2X1 U1862 (.Y(n1393), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN563_n667), 
	.A1N(key_mem[899]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1863 (.Y(n1392), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN562_n666), 
	.A1N(key_mem[900]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1864 (.Y(n1391), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN566_n665), 
	.A1N(key_mem[901]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1865 (.Y(n1390), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN572_n664), 
	.A1N(key_mem[902]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1866 (.Y(n1389), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN324_n663), 
	.A1N(key_mem[903]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1867 (.Y(n1388), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN325_n662), 
	.A1N(key_mem[904]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1868 (.Y(n1387), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN323_n661), 
	.A1N(key_mem[905]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1869 (.Y(n1386), 
	.B1(n676), 
	.B0(FE_PHN541_n660), 
	.A1N(key_mem[906]), 
	.A0N(n676));
   OAI2BB2X1 U1870 (.Y(n1385), 
	.B1(n676), 
	.B0(FE_PHN554_n659), 
	.A1N(key_mem[907]), 
	.A0N(n676));
   OAI2BB2X1 U1871 (.Y(n1384), 
	.B1(n676), 
	.B0(FE_PHN560_n658), 
	.A1N(key_mem[908]), 
	.A0N(n676));
   OAI2BB2X1 U1872 (.Y(n1383), 
	.B1(n676), 
	.B0(FE_PHN552_n657), 
	.A1N(key_mem[909]), 
	.A0N(n676));
   OAI2BB2X1 U1873 (.Y(n1380), 
	.B1(FE_OFN76_n676), 
	.B0(FE_PHN573_n654), 
	.A1N(key_mem[912]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U1874 (.Y(n1376), 
	.B1(FE_OFN76_n676), 
	.B0(FE_PHN579_n650), 
	.A1N(key_mem[916]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U1875 (.Y(n1364), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN383_n638), 
	.A1N(key_mem[928]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1876 (.Y(n1363), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN380_n637), 
	.A1N(key_mem[929]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1877 (.Y(n1362), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN381_n636), 
	.A1N(key_mem[930]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1878 (.Y(n1361), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN379_n635), 
	.A1N(key_mem[931]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1879 (.Y(n1360), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN394_n634), 
	.A1N(key_mem[932]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1880 (.Y(n1359), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN391_n633), 
	.A1N(key_mem[933]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1881 (.Y(n1358), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN396_n632), 
	.A1N(key_mem[934]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1882 (.Y(n1357), 
	.B1(FE_OFN77_n676), 
	.B0(n631), 
	.A1N(key_mem[935]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1883 (.Y(n1356), 
	.B1(FE_OFN77_n676), 
	.B0(n630), 
	.A1N(key_mem[936]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1884 (.Y(n1355), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN705_n629), 
	.A1N(key_mem[937]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1885 (.Y(n1354), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN390_n628), 
	.A1N(key_mem[938]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1886 (.Y(n1353), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN398_n627), 
	.A1N(key_mem[939]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1887 (.Y(n1352), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN388_n626), 
	.A1N(key_mem[940]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1888 (.Y(n1351), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN387_n625), 
	.A1N(key_mem[941]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1889 (.Y(n1350), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN409_n624), 
	.A1N(key_mem[942]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1890 (.Y(n1349), 
	.B1(FE_OFN77_n676), 
	.B0(n623), 
	.A1N(key_mem[943]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1891 (.Y(n1348), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN403_n622), 
	.A1N(key_mem[944]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1892 (.Y(n1347), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN402_n621), 
	.A1N(key_mem[945]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1893 (.Y(n1346), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN384_n620), 
	.A1N(key_mem[946]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1894 (.Y(n1345), 
	.B1(n676), 
	.B0(FE_PHN382_n619), 
	.A1N(key_mem[947]), 
	.A0N(n676));
   OAI2BB2X1 U1895 (.Y(n1343), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN385_n617), 
	.A1N(key_mem[949]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1896 (.Y(n1342), 
	.B1(FE_OFN77_n676), 
	.B0(n616), 
	.A1N(key_mem[950]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1897 (.Y(n1341), 
	.B1(FE_OFN77_n676), 
	.B0(n615), 
	.A1N(key_mem[951]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1898 (.Y(n1332), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN540_n606), 
	.A1N(key_mem[960]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1899 (.Y(n1331), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN555_n605), 
	.A1N(key_mem[961]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1900 (.Y(n1330), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN538_n604), 
	.A1N(key_mem[962]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1901 (.Y(n1329), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN546_n603), 
	.A1N(key_mem[963]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1902 (.Y(n1328), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN557_n602), 
	.A1N(key_mem[964]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1903 (.Y(n1327), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN561_n601), 
	.A1N(key_mem[965]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1904 (.Y(n1325), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN545_n599), 
	.A1N(key_mem[967]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1905 (.Y(n1324), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN559_n598), 
	.A1N(key_mem[968]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1906 (.Y(n1323), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN416_n597), 
	.A1N(FE_PHN3433_key_mem_969_), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1907 (.Y(n1322), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN565_n596), 
	.A1N(key_mem[970]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1908 (.Y(n1321), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN556_n595), 
	.A1N(key_mem[971]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1909 (.Y(n1320), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN575_n594), 
	.A1N(key_mem[972]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1910 (.Y(n1319), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN577_n593), 
	.A1N(key_mem[973]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1911 (.Y(n1318), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN420_n592), 
	.A1N(key_mem[974]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1912 (.Y(n1317), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN417_n591), 
	.A1N(key_mem[975]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1913 (.Y(n1314), 
	.B1(n676), 
	.B0(FE_PHN543_n588), 
	.A1N(key_mem[978]), 
	.A0N(n676));
   OAI2BB2X1 U1914 (.Y(n1313), 
	.B1(n676), 
	.B0(FE_PHN549_n587), 
	.A1N(key_mem[979]), 
	.A0N(n676));
   OAI2BB2X1 U1915 (.Y(n1311), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN539_n585), 
	.A1N(key_mem[981]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1916 (.Y(n1310), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN576_n584), 
	.A1N(key_mem[982]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U1917 (.Y(n1309), 
	.B1(n676), 
	.B0(FE_PHN574_n583), 
	.A1N(key_mem[983]), 
	.A0N(n676));
   OAI2BB2X1 U1918 (.Y(n1300), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN609_n574), 
	.A1N(key_mem[992]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1919 (.Y(n1297), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN606_n571), 
	.A1N(key_mem[995]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1920 (.Y(n1292), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN607_n566), 
	.A1N(key_mem[1000]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U1921 (.Y(n1291), 
	.B1(n676), 
	.B0(n565), 
	.A1N(key_mem[1001]), 
	.A0N(n676));
   OAI2BB2X1 U1922 (.Y(n1290), 
	.B1(n676), 
	.B0(FE_PHN608_n564), 
	.A1N(FE_PHN3426_key_mem_1002_), 
	.A0N(n676));
   OAI2BB2X1 U1923 (.Y(n1289), 
	.B1(n676), 
	.B0(FE_PHN615_n563), 
	.A1N(key_mem[1003]), 
	.A0N(n676));
   OAI2BB2X1 U1924 (.Y(n1287), 
	.B1(n676), 
	.B0(FE_PHN621_n561), 
	.A1N(key_mem[1005]), 
	.A0N(n676));
   OAI2BB2X1 U1925 (.Y(n1285), 
	.B1(FE_OFN76_n676), 
	.B0(n559), 
	.A1N(FE_PHN3431_key_mem_1007_), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U1926 (.Y(n1012), 
	.B1(FE_OFN88_n1), 
	.B0(FE_PHN553_n670), 
	.A1N(key_mem[1280]), 
	.A0N(FE_OFN88_n1));
   OAI2BB2X1 U1927 (.Y(n1011), 
	.B1(FE_OFN86_n1), 
	.B0(FE_PHN537_n669), 
	.A1N(key_mem[1281]), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U1928 (.Y(n1010), 
	.B1(n1), 
	.B0(FE_PHN550_n668), 
	.A1N(FE_PHN2825_key_mem_1282_), 
	.A0N(n1));
   OAI2BB2X1 U1929 (.Y(n1009), 
	.B1(FE_OFN89_n1), 
	.B0(FE_PHN563_n667), 
	.A1N(key_mem[1283]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U1930 (.Y(n1008), 
	.B1(FE_OFN89_n1), 
	.B0(FE_PHN562_n666), 
	.A1N(key_mem[1284]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U1931 (.Y(n1007), 
	.B1(FE_OFN87_n1), 
	.B0(FE_PHN566_n665), 
	.A1N(key_mem[1285]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U1932 (.Y(n1006), 
	.B1(FE_OFN86_n1), 
	.B0(FE_PHN572_n664), 
	.A1N(key_mem[1286]), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U1933 (.Y(n1005), 
	.B1(FE_OFN88_n1), 
	.B0(FE_PHN324_n663), 
	.A1N(key_mem[1287]), 
	.A0N(FE_OFN88_n1));
   OAI2BB2X1 U1934 (.Y(n1004), 
	.B1(FE_OFN86_n1), 
	.B0(FE_PHN325_n662), 
	.A1N(key_mem[1288]), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U1935 (.Y(n1003), 
	.B1(FE_OFN86_n1), 
	.B0(FE_PHN323_n661), 
	.A1N(FE_PHN3205_key_mem_1289_), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U1936 (.Y(n1002), 
	.B1(n1), 
	.B0(FE_PHN541_n660), 
	.A1N(FE_PHN3285_key_mem_1290_), 
	.A0N(n1));
   OAI2BB2X1 U1937 (.Y(n1001), 
	.B1(n1), 
	.B0(FE_PHN554_n659), 
	.A1N(key_mem[1291]), 
	.A0N(n1));
   OAI2BB2X1 U1938 (.Y(n1000), 
	.B1(n1), 
	.B0(FE_PHN560_n658), 
	.A1N(key_mem[1292]), 
	.A0N(n1));
   OAI2BB2X1 U1939 (.Y(n999), 
	.B1(n1), 
	.B0(FE_PHN552_n657), 
	.A1N(key_mem[1293]), 
	.A0N(n1));
   OAI2BB2X1 U1940 (.Y(n996), 
	.B1(FE_OFN85_n1), 
	.B0(FE_PHN573_n654), 
	.A1N(key_mem[1296]), 
	.A0N(FE_OFN85_n1));
   OAI2BB2X1 U1941 (.Y(n992), 
	.B1(FE_OFN85_n1), 
	.B0(FE_PHN579_n650), 
	.A1N(key_mem[1300]), 
	.A0N(FE_OFN85_n1));
   OAI2BB2X1 U1942 (.Y(n980), 
	.B1(FE_OFN86_n1), 
	.B0(FE_PHN383_n638), 
	.A1N(key_mem[1312]), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U1943 (.Y(n979), 
	.B1(FE_OFN86_n1), 
	.B0(FE_PHN380_n637), 
	.A1N(key_mem[1313]), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U1944 (.Y(n978), 
	.B1(FE_OFN88_n1), 
	.B0(FE_PHN381_n636), 
	.A1N(key_mem[1314]), 
	.A0N(FE_OFN88_n1));
   OAI2BB2X1 U1945 (.Y(n977), 
	.B1(FE_OFN86_n1), 
	.B0(FE_PHN379_n635), 
	.A1N(key_mem[1315]), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U1946 (.Y(n976), 
	.B1(FE_OFN86_n1), 
	.B0(FE_PHN394_n634), 
	.A1N(key_mem[1316]), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U1947 (.Y(n975), 
	.B1(FE_OFN88_n1), 
	.B0(FE_PHN391_n633), 
	.A1N(key_mem[1317]), 
	.A0N(FE_OFN88_n1));
   OAI2BB2X1 U1949 (.Y(n974), 
	.B1(FE_OFN86_n1), 
	.B0(FE_PHN396_n632), 
	.A1N(key_mem[1318]), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U1950 (.Y(n973), 
	.B1(FE_OFN89_n1), 
	.B0(n631), 
	.A1N(key_mem[1319]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U1951 (.Y(n972), 
	.B1(FE_OFN89_n1), 
	.B0(n630), 
	.A1N(key_mem[1320]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U1952 (.Y(n971), 
	.B1(FE_OFN89_n1), 
	.B0(FE_PHN705_n629), 
	.A1N(key_mem[1321]), 
	.A0N(FE_OFN88_n1));
   OAI2BB2X1 U1953 (.Y(n970), 
	.B1(FE_OFN89_n1), 
	.B0(FE_PHN390_n628), 
	.A1N(key_mem[1322]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U1954 (.Y(n969), 
	.B1(FE_OFN87_n1), 
	.B0(FE_PHN398_n627), 
	.A1N(key_mem[1323]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U1955 (.Y(n968), 
	.B1(FE_OFN89_n1), 
	.B0(FE_PHN388_n626), 
	.A1N(key_mem[1324]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U1956 (.Y(n967), 
	.B1(FE_OFN89_n1), 
	.B0(FE_PHN387_n625), 
	.A1N(key_mem[1325]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U1957 (.Y(n966), 
	.B1(FE_OFN89_n1), 
	.B0(FE_PHN409_n624), 
	.A1N(key_mem[1326]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U1958 (.Y(n965), 
	.B1(FE_OFN89_n1), 
	.B0(n623), 
	.A1N(key_mem[1327]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U1959 (.Y(n964), 
	.B1(FE_OFN89_n1), 
	.B0(FE_PHN403_n622), 
	.A1N(key_mem[1328]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U1960 (.Y(n963), 
	.B1(FE_OFN89_n1), 
	.B0(FE_PHN402_n621), 
	.A1N(key_mem[1329]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U1961 (.Y(n962), 
	.B1(FE_OFN89_n1), 
	.B0(FE_PHN384_n620), 
	.A1N(key_mem[1330]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U1962 (.Y(n961), 
	.B1(FE_OFN87_n1), 
	.B0(FE_PHN382_n619), 
	.A1N(key_mem[1331]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U1963 (.Y(n959), 
	.B1(FE_OFN87_n1), 
	.B0(FE_PHN385_n617), 
	.A1N(key_mem[1333]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U1964 (.Y(n958), 
	.B1(FE_OFN87_n1), 
	.B0(n616), 
	.A1N(key_mem[1334]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U1965 (.Y(n957), 
	.B1(FE_OFN87_n1), 
	.B0(n615), 
	.A1N(key_mem[1335]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U1966 (.Y(n948), 
	.B1(FE_OFN88_n1), 
	.B0(FE_PHN540_n606), 
	.A1N(FE_PHN969_key_mem_1344_), 
	.A0N(FE_OFN88_n1));
   OAI2BB2X1 U1967 (.Y(n947), 
	.B1(FE_OFN88_n1), 
	.B0(FE_PHN555_n605), 
	.A1N(FE_PHN774_key_mem_1345_), 
	.A0N(FE_OFN88_n1));
   OAI2BB2X1 U1968 (.Y(n946), 
	.B1(FE_OFN88_n1), 
	.B0(FE_PHN538_n604), 
	.A1N(key_mem[1346]), 
	.A0N(FE_OFN88_n1));
   OAI2BB2X1 U1969 (.Y(n945), 
	.B1(FE_OFN88_n1), 
	.B0(FE_PHN546_n603), 
	.A1N(key_mem[1347]), 
	.A0N(FE_OFN88_n1));
   OAI2BB2X1 U1970 (.Y(n944), 
	.B1(FE_OFN88_n1), 
	.B0(FE_PHN557_n602), 
	.A1N(key_mem[1348]), 
	.A0N(FE_OFN88_n1));
   OAI2BB2X1 U1971 (.Y(n943), 
	.B1(FE_OFN89_n1), 
	.B0(FE_PHN561_n601), 
	.A1N(key_mem[1349]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U1972 (.Y(n941), 
	.B1(FE_OFN88_n1), 
	.B0(FE_PHN545_n599), 
	.A1N(FE_PHN2828_key_mem_1351_), 
	.A0N(FE_OFN88_n1));
   OAI2BB2X1 U1973 (.Y(n940), 
	.B1(FE_OFN88_n1), 
	.B0(FE_PHN559_n598), 
	.A1N(key_mem[1352]), 
	.A0N(FE_OFN88_n1));
   OAI2BB2X1 U1974 (.Y(n939), 
	.B1(FE_OFN86_n1), 
	.B0(FE_PHN416_n597), 
	.A1N(FE_PHN2841_key_mem_1353_), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U1975 (.Y(n938), 
	.B1(FE_OFN86_n1), 
	.B0(FE_PHN565_n596), 
	.A1N(key_mem[1354]), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U1976 (.Y(n937), 
	.B1(FE_OFN86_n1), 
	.B0(FE_PHN556_n595), 
	.A1N(key_mem[1355]), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U1977 (.Y(n936), 
	.B1(FE_OFN86_n1), 
	.B0(FE_PHN575_n594), 
	.A1N(key_mem[1356]), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U1978 (.Y(n935), 
	.B1(FE_OFN86_n1), 
	.B0(FE_PHN577_n593), 
	.A1N(key_mem[1357]), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U1979 (.Y(n934), 
	.B1(FE_OFN88_n1), 
	.B0(FE_PHN420_n592), 
	.A1N(key_mem[1358]), 
	.A0N(FE_OFN88_n1));
   OAI2BB2X1 U1980 (.Y(n933), 
	.B1(n2624), 
	.B0(FE_PHN417_n591), 
	.A1N(key_mem[1359]), 
	.A0N(FE_OFN88_n1));
   OAI2BB2X1 U1981 (.Y(n930), 
	.B1(n2624), 
	.B0(FE_PHN543_n588), 
	.A1N(key_mem[1362]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U1982 (.Y(n929), 
	.B1(n2624), 
	.B0(FE_PHN549_n587), 
	.A1N(key_mem[1363]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U1983 (.Y(n927), 
	.B1(n2624), 
	.B0(FE_PHN539_n585), 
	.A1N(key_mem[1365]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U1984 (.Y(n926), 
	.B1(n2624), 
	.B0(FE_PHN576_n584), 
	.A1N(key_mem[1366]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U1985 (.Y(n925), 
	.B1(n2624), 
	.B0(FE_PHN574_n583), 
	.A1N(key_mem[1367]), 
	.A0N(n1));
   OAI2BB2X1 U1986 (.Y(n916), 
	.B1(n2623), 
	.B0(FE_PHN609_n574), 
	.A1N(key_mem[1376]), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U1987 (.Y(n913), 
	.B1(n2623), 
	.B0(FE_PHN606_n571), 
	.A1N(FE_PHN932_key_mem_1379_), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U1988 (.Y(n908), 
	.B1(n2622), 
	.B0(FE_PHN607_n566), 
	.A1N(key_mem[1384]), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U1989 (.Y(n907), 
	.B1(n2622), 
	.B0(n565), 
	.A1N(key_mem[1385]), 
	.A0N(n1));
   OAI2BB2X1 U1990 (.Y(n906), 
	.B1(n2622), 
	.B0(FE_PHN608_n564), 
	.A1N(FE_PHN2810_key_mem_1386_), 
	.A0N(n1));
   OAI2BB2X1 U1991 (.Y(n905), 
	.B1(n2622), 
	.B0(FE_PHN615_n563), 
	.A1N(key_mem[1387]), 
	.A0N(n1));
   OAI2BB2X1 U1992 (.Y(n903), 
	.B1(n2622), 
	.B0(FE_PHN621_n561), 
	.A1N(key_mem[1389]), 
	.A0N(n1));
   OAI2BB2X1 U1993 (.Y(n901), 
	.B1(n2622), 
	.B0(n559), 
	.A1N(FE_PHN3419_key_mem_1391_), 
	.A0N(FE_OFN85_n1));
   AOI22X1 U1995 (.Y(n573), 
	.B1(n2652), 
	.B0(key[97]), 
	.A1(n729), 
	.A0(FE_OFN91_n690));
   AOI22X1 U1997 (.Y(n572), 
	.B1(n2651), 
	.B0(key[98]), 
	.A1(n728), 
	.A0(FE_OFN90_n690));
   AOI22X1 U1999 (.Y(n571), 
	.B1(n2651), 
	.B0(key[99]), 
	.A1(n727), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2001 (.Y(n570), 
	.B1(n2650), 
	.B0(key[100]), 
	.A1(n726), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2003 (.Y(n569), 
	.B1(n2650), 
	.B0(key[101]), 
	.A1(n725), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2005 (.Y(n567), 
	.B1(n2649), 
	.B0(key[103]), 
	.A1(n723), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2007 (.Y(n566), 
	.B1(n2648), 
	.B0(key[104]), 
	.A1(n722), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2009 (.Y(n565), 
	.B1(n2648), 
	.B0(key[105]), 
	.A1(n721), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2011 (.Y(n564), 
	.B1(n2647), 
	.B0(key[106]), 
	.A1(n720), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2013 (.Y(n563), 
	.B1(n2647), 
	.B0(key[107]), 
	.A1(n719), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2015 (.Y(n562), 
	.B1(n2646), 
	.B0(key[108]), 
	.A1(n718), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2017 (.Y(n561), 
	.B1(n2646), 
	.B0(key[109]), 
	.A1(n717), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2019 (.Y(n560), 
	.B1(n2645), 
	.B0(key[110]), 
	.A1(n716), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2021 (.Y(n559), 
	.B1(n2645), 
	.B0(key[111]), 
	.A1(n715), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2023 (.Y(n556), 
	.B1(n2643), 
	.B0(key[114]), 
	.A1(n712), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2025 (.Y(n555), 
	.B1(n2643), 
	.B0(key[115]), 
	.A1(n711), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2027 (.Y(n553), 
	.B1(n2642), 
	.B0(key[117]), 
	.A1(n709), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2029 (.Y(n552), 
	.B1(n2641), 
	.B0(key[118]), 
	.A1(n708), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2031 (.Y(n551), 
	.B1(n2641), 
	.B0(key[119]), 
	.A1(n707), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2033 (.Y(n575), 
	.B1(n2653), 
	.B0(key[95]), 
	.A1(n731), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2035 (.Y(n582), 
	.B1(n2656), 
	.B0(key[88]), 
	.A1(n738), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2037 (.Y(n576), 
	.B1(n2653), 
	.B0(key[94]), 
	.A1(n732), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2039 (.Y(n577), 
	.B1(n2654), 
	.B0(key[93]), 
	.A1(n733), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2041 (.Y(n578), 
	.B1(n2654), 
	.B0(key[92]), 
	.A1(n734), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2043 (.Y(n579), 
	.B1(n2655), 
	.B0(key[91]), 
	.A1(n735), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2045 (.Y(n581), 
	.B1(n2656), 
	.B0(key[89]), 
	.A1(n737), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2047 (.Y(n638), 
	.B1(n2684), 
	.B0(key[32]), 
	.A1(n810), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2049 (.Y(n637), 
	.B1(n2684), 
	.B0(key[33]), 
	.A1(n809), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2051 (.Y(n636), 
	.B1(n2683), 
	.B0(key[34]), 
	.A1(n808), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2053 (.Y(n635), 
	.B1(n2683), 
	.B0(key[35]), 
	.A1(n807), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2055 (.Y(n634), 
	.B1(n2682), 
	.B0(key[36]), 
	.A1(n806), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2057 (.Y(n633), 
	.B1(n2682), 
	.B0(key[37]), 
	.A1(n805), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2059 (.Y(n632), 
	.B1(n2681), 
	.B0(key[38]), 
	.A1(n804), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2061 (.Y(n631), 
	.B1(n2681), 
	.B0(key[39]), 
	.A1(n803), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2063 (.Y(n630), 
	.B1(n2680), 
	.B0(key[40]), 
	.A1(n802), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2065 (.Y(n629), 
	.B1(n2680), 
	.B0(key[41]), 
	.A1(n801), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2067 (.Y(n628), 
	.B1(n2679), 
	.B0(key[42]), 
	.A1(n800), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2069 (.Y(n627), 
	.B1(n2679), 
	.B0(key[43]), 
	.A1(n799), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2071 (.Y(n626), 
	.B1(n2678), 
	.B0(key[44]), 
	.A1(n798), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2073 (.Y(n625), 
	.B1(n2678), 
	.B0(key[45]), 
	.A1(n797), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2075 (.Y(n624), 
	.B1(n2677), 
	.B0(key[46]), 
	.A1(n796), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2077 (.Y(n623), 
	.B1(n2677), 
	.B0(key[47]), 
	.A1(n795), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2080 (.Y(n622), 
	.B1(n2676), 
	.B0(key[48]), 
	.A1(n794), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2082 (.Y(n621), 
	.B1(n2676), 
	.B0(key[49]), 
	.A1(n793), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2084 (.Y(n620), 
	.B1(n2675), 
	.B0(key[50]), 
	.A1(n792), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2086 (.Y(n619), 
	.B1(n2675), 
	.B0(key[51]), 
	.A1(n791), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2088 (.Y(n618), 
	.B1(n2674), 
	.B0(key[52]), 
	.A1(n790), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2090 (.Y(n617), 
	.B1(n2674), 
	.B0(key[53]), 
	.A1(n789), 
	.A0(FE_OFN90_n690));
   AOI22X1 U2092 (.Y(n616), 
	.B1(n2673), 
	.B0(key[54]), 
	.A1(n788), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2094 (.Y(n615), 
	.B1(n2673), 
	.B0(key[55]), 
	.A1(n787), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2096 (.Y(n543), 
	.B1(n691), 
	.B0(FE_OFN91_n690), 
	.A1(n2637), 
	.A0(key[127]));
   XOR2X1 U2097 (.Y(n691), 
	.B(n692), 
	.A(FE_PHN1434_prev_key1_reg_127_));
   AOI22X1 U2099 (.Y(n640), 
	.B1(n2685), 
	.B0(key[30]), 
	.A1(n813), 
	.A0(FE_OFN91_n690));
   XNOR2X1 U2100 (.Y(n813), 
	.B(n732), 
	.A(n814));
   XNOR2X1 U2101 (.Y(n814), 
	.B(sboxw[30]), 
	.A(FE_PHN740_prev_key1_reg_62_));
   AOI22X1 U2103 (.Y(n608), 
	.B1(n2669), 
	.B0(key[62]), 
	.A1(n766), 
	.A0(FE_OFN91_n690));
   XNOR2X1 U2104 (.Y(n766), 
	.B(n768), 
	.A(n767));
   XNOR2X1 U2105 (.Y(n767), 
	.B(n694), 
	.A(FE_PHN740_prev_key1_reg_62_));
   AOI22X1 U2107 (.Y(n610), 
	.B1(n2670), 
	.B0(key[60]), 
	.A1(n772), 
	.A0(FE_OFN90_n690));
   XNOR2X1 U2108 (.Y(n772), 
	.B(n774), 
	.A(n773));
   XNOR2X1 U2109 (.Y(n773), 
	.B(n698), 
	.A(FE_PHN741_prev_key1_reg_60_));
   AOI22X1 U2111 (.Y(n546), 
	.B1(n697), 
	.B0(FE_OFN90_n690), 
	.A1(n2638), 
	.A0(key[124]));
   XOR2X1 U2112 (.Y(n697), 
	.B(n698), 
	.A(FE_PHN1421_prev_key1_reg_124_));
   AOI22X1 U2114 (.Y(n548), 
	.B1(n701), 
	.B0(FE_OFN90_n690), 
	.A1(n2639), 
	.A0(key[122]));
   XOR2X1 U2115 (.Y(n701), 
	.B(n702), 
	.A(FE_PHN1392_prev_key1_reg_122_));
   AOI22X1 U2117 (.Y(n666), 
	.B1(n2698), 
	.B0(key[4]), 
	.A1(n865), 
	.A0(FE_OFN90_n690));
   XOR2X1 U2118 (.Y(n865), 
	.B(n806), 
	.A(FE_PHN2003_keymem_sboxw_4_));
   AOI22X1 U2120 (.Y(n665), 
	.B1(n2698), 
	.B0(key[5]), 
	.A1(n863), 
	.A0(FE_OFN90_n690));
   XOR2X1 U2121 (.Y(n863), 
	.B(n805), 
	.A(FE_PHN2006_keymem_sboxw_5_));
   AOI22X1 U2123 (.Y(n664), 
	.B1(n2697), 
	.B0(key[6]), 
	.A1(n861), 
	.A0(FE_OFN91_n690));
   XOR2X1 U2124 (.Y(n861), 
	.B(n804), 
	.A(sboxw[6]));
   AOI22X1 U2126 (.Y(n663), 
	.B1(n2697), 
	.B0(key[7]), 
	.A1(n859), 
	.A0(FE_OFN91_n690));
   XOR2X1 U2127 (.Y(n859), 
	.B(n803), 
	.A(sboxw[7]));
   AOI22X1 U2129 (.Y(n656), 
	.B1(n2693), 
	.B0(key[14]), 
	.A1(n845), 
	.A0(FE_OFN91_n690));
   XOR2X1 U2130 (.Y(n845), 
	.B(n796), 
	.A(sboxw[14]));
   AOI22X1 U2132 (.Y(n654), 
	.B1(n2692), 
	.B0(key[16]), 
	.A1(n841), 
	.A0(FE_OFN91_n690));
   XOR2X1 U2133 (.Y(n841), 
	.B(n794), 
	.A(sboxw[16]));
   AOI22X1 U2135 (.Y(n653), 
	.B1(n2692), 
	.B0(key[17]), 
	.A1(n839), 
	.A0(FE_OFN91_n690));
   XOR2X1 U2136 (.Y(n839), 
	.B(n793), 
	.A(FE_PHN1998_keymem_sboxw_17_));
   AOI22X1 U2138 (.Y(n652), 
	.B1(n2691), 
	.B0(key[18]), 
	.A1(n837), 
	.A0(FE_OFN90_n690));
   XOR2X1 U2139 (.Y(n837), 
	.B(n792), 
	.A(FE_PHN1958_keymem_sboxw_18_));
   AOI22X1 U2141 (.Y(n651), 
	.B1(n2691), 
	.B0(key[19]), 
	.A1(n835), 
	.A0(FE_OFN90_n690));
   XOR2X1 U2142 (.Y(n835), 
	.B(n791), 
	.A(sboxw[19]));
   AOI22X1 U2144 (.Y(n650), 
	.B1(n2690), 
	.B0(key[20]), 
	.A1(n833), 
	.A0(FE_OFN90_n690));
   XOR2X1 U2145 (.Y(n833), 
	.B(n790), 
	.A(FE_PHN2005_keymem_sboxw_20_));
   AOI22X1 U2147 (.Y(n649), 
	.B1(n2690), 
	.B0(key[21]), 
	.A1(n831), 
	.A0(FE_OFN90_n690));
   XOR2X1 U2148 (.Y(n831), 
	.B(n789), 
	.A(sboxw[21]));
   AOI22X1 U2150 (.Y(n648), 
	.B1(n2689), 
	.B0(key[22]), 
	.A1(n829), 
	.A0(FE_OFN91_n690));
   XOR2X1 U2151 (.Y(n829), 
	.B(n788), 
	.A(FE_PHN1965_keymem_sboxw_22_));
   AOI22X1 U2153 (.Y(n647), 
	.B1(n2689), 
	.B0(key[23]), 
	.A1(n827), 
	.A0(FE_OFN91_n690));
   XOR2X1 U2154 (.Y(n827), 
	.B(n787), 
	.A(sboxw[23]));
   AOI22X1 U2156 (.Y(n606), 
	.B1(n2668), 
	.B0(key[64]), 
	.A1(n762), 
	.A0(FE_OFN91_n690));
   XOR2X1 U2157 (.Y(n762), 
	.B(n730), 
	.A(FE_PHN1441_prev_key1_reg_64_));
   AOI22X1 U2159 (.Y(n605), 
	.B1(n2668), 
	.B0(key[65]), 
	.A1(n761), 
	.A0(FE_OFN91_n690));
   XOR2X1 U2160 (.Y(n761), 
	.B(n729), 
	.A(FE_PHN1394_prev_key1_reg_65_));
   AOI22X1 U2162 (.Y(n604), 
	.B1(n2667), 
	.B0(key[66]), 
	.A1(n760), 
	.A0(FE_OFN90_n690));
   XOR2X1 U2163 (.Y(n760), 
	.B(n728), 
	.A(FE_PHN1442_prev_key1_reg_66_));
   AOI22X1 U2165 (.Y(n603), 
	.B1(n2667), 
	.B0(key[67]), 
	.A1(n759), 
	.A0(FE_OFN90_n690));
   XOR2X1 U2166 (.Y(n759), 
	.B(n727), 
	.A(FE_PHN1444_prev_key1_reg_67_));
   AOI22X1 U2168 (.Y(n602), 
	.B1(n2666), 
	.B0(key[68]), 
	.A1(n758), 
	.A0(FE_OFN90_n690));
   XOR2X1 U2169 (.Y(n758), 
	.B(n726), 
	.A(FE_PHN1446_prev_key1_reg_68_));
   AOI22X1 U2171 (.Y(n601), 
	.B1(n2666), 
	.B0(key[69]), 
	.A1(n757), 
	.A0(FE_OFN90_n690));
   XOR2X1 U2172 (.Y(n757), 
	.B(n725), 
	.A(FE_PHN1445_prev_key1_reg_69_));
   AOI22X1 U2174 (.Y(n600), 
	.B1(n2665), 
	.B0(key[70]), 
	.A1(n756), 
	.A0(FE_OFN91_n690));
   XOR2X1 U2175 (.Y(n756), 
	.B(n724), 
	.A(prev_key1_reg[70]));
   AOI22X1 U2177 (.Y(n599), 
	.B1(n2665), 
	.B0(key[71]), 
	.A1(n755), 
	.A0(FE_OFN91_n690));
   XOR2X1 U2178 (.Y(n755), 
	.B(n723), 
	.A(FE_PHN1406_prev_key1_reg_71_));
   AOI22X1 U2180 (.Y(n598), 
	.B1(n2664), 
	.B0(key[72]), 
	.A1(n754), 
	.A0(FE_OFN91_n690));
   XOR2X1 U2181 (.Y(n754), 
	.B(n722), 
	.A(FE_PHN1404_prev_key1_reg_72_));
   AOI22X1 U2183 (.Y(n597), 
	.B1(n2664), 
	.B0(key[73]), 
	.A1(n753), 
	.A0(FE_OFN91_n690));
   XOR2X1 U2184 (.Y(n753), 
	.B(n721), 
	.A(FE_PHN1401_prev_key1_reg_73_));
   AOI22X1 U2186 (.Y(n596), 
	.B1(n2663), 
	.B0(key[74]), 
	.A1(n752), 
	.A0(FE_OFN90_n690));
   XOR2X1 U2187 (.Y(n752), 
	.B(n720), 
	.A(FE_PHN1408_prev_key1_reg_74_));
   AOI22X1 U2189 (.Y(n595), 
	.B1(n2663), 
	.B0(key[75]), 
	.A1(n751), 
	.A0(FE_OFN90_n690));
   XOR2X1 U2190 (.Y(n751), 
	.B(n719), 
	.A(FE_PHN1415_prev_key1_reg_75_));
   AOI22X1 U2192 (.Y(n594), 
	.B1(n2662), 
	.B0(key[76]), 
	.A1(n750), 
	.A0(FE_OFN90_n690));
   XOR2X1 U2193 (.Y(n750), 
	.B(n718), 
	.A(FE_PHN1429_prev_key1_reg_76_));
   AOI22X1 U2195 (.Y(n593), 
	.B1(n2662), 
	.B0(key[77]), 
	.A1(n749), 
	.A0(FE_OFN90_n690));
   XOR2X1 U2196 (.Y(n749), 
	.B(n717), 
	.A(FE_PHN1397_prev_key1_reg_77_));
   AOI22X1 U2198 (.Y(n592), 
	.B1(n2661), 
	.B0(key[78]), 
	.A1(n748), 
	.A0(FE_OFN91_n690));
   XOR2X1 U2199 (.Y(n748), 
	.B(n716), 
	.A(FE_PHN1402_prev_key1_reg_78_));
   AOI22X1 U2201 (.Y(n591), 
	.B1(n2661), 
	.B0(key[79]), 
	.A1(n747), 
	.A0(FE_OFN91_n690));
   XOR2X1 U2202 (.Y(n747), 
	.B(n715), 
	.A(FE_PHN1393_prev_key1_reg_79_));
   AOI22X1 U2204 (.Y(n590), 
	.B1(n2660), 
	.B0(key[80]), 
	.A1(n746), 
	.A0(FE_OFN91_n690));
   XOR2X1 U2205 (.Y(n746), 
	.B(n714), 
	.A(FE_PHN1414_prev_key1_reg_80_));
   AOI22X1 U2207 (.Y(n589), 
	.B1(n2660), 
	.B0(key[81]), 
	.A1(n745), 
	.A0(FE_OFN91_n690));
   XOR2X1 U2208 (.Y(n745), 
	.B(n713), 
	.A(FE_PHN1425_prev_key1_reg_81_));
   AOI22X1 U2210 (.Y(n588), 
	.B1(n2659), 
	.B0(key[82]), 
	.A1(n744), 
	.A0(FE_OFN90_n690));
   XOR2X1 U2211 (.Y(n744), 
	.B(n712), 
	.A(FE_PHN1405_prev_key1_reg_82_));
   AOI22X1 U2213 (.Y(n587), 
	.B1(n2659), 
	.B0(key[83]), 
	.A1(n743), 
	.A0(FE_OFN90_n690));
   XOR2X1 U2214 (.Y(n743), 
	.B(n711), 
	.A(FE_PHN1388_prev_key1_reg_83_));
   AOI22X1 U2216 (.Y(n586), 
	.B1(n2658), 
	.B0(key[84]), 
	.A1(n742), 
	.A0(FE_OFN90_n690));
   XOR2X1 U2217 (.Y(n742), 
	.B(n710), 
	.A(FE_PHN1375_prev_key1_reg_84_));
   AOI22X1 U2219 (.Y(n585), 
	.B1(n2658), 
	.B0(key[85]), 
	.A1(n741), 
	.A0(FE_OFN90_n690));
   XOR2X1 U2220 (.Y(n741), 
	.B(n709), 
	.A(FE_PHN1412_prev_key1_reg_85_));
   AOI22X1 U2222 (.Y(n584), 
	.B1(n2657), 
	.B0(key[86]), 
	.A1(n740), 
	.A0(FE_OFN91_n690));
   XOR2X1 U2223 (.Y(n740), 
	.B(n708), 
	.A(FE_PHN360_prev_key1_reg_86_));
   AOI22X1 U2225 (.Y(n583), 
	.B1(n2657), 
	.B0(key[87]), 
	.A1(n739), 
	.A0(FE_OFN91_n690));
   XOR2X1 U2226 (.Y(n739), 
	.B(n707), 
	.A(FE_PHN359_prev_key1_reg_87_));
   OAI2BB2X1 U2227 (.Y(n1216), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN389_n618), 
	.A1N(FE_PHN1798_key_mem_1076_), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U2228 (.Y(n1198), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN578_n600), 
	.A1N(FE_PHN1863_key_mem_1094_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U2229 (.Y(n1188), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN421_n590), 
	.A1N(FE_PHN1821_key_mem_1104_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U2230 (.Y(n1187), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN419_n589), 
	.A1N(FE_PHN1745_key_mem_1105_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U2231 (.Y(n1184), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN542_n586), 
	.A1N(key_mem[1108]), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U2232 (.Y(n1171), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN610_n573), 
	.A1N(FE_PHN1850_key_mem_1121_), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U2233 (.Y(n1170), 
	.B1(FE_OFN96_n674), 
	.B0(FE_PHN612_n572), 
	.A1N(key_mem[1122]), 
	.A0N(FE_OFN96_n674));
   OAI2BB2X1 U2234 (.Y(n1168), 
	.B1(n674), 
	.B0(FE_PHN617_n570), 
	.A1N(key_mem[1124]), 
	.A0N(n674));
   OAI2BB2X1 U2235 (.Y(n1167), 
	.B1(n674), 
	.B0(FE_PHN613_n569), 
	.A1N(key_mem[1125]), 
	.A0N(n674));
   OAI2BB2X1 U2236 (.Y(n1166), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN605_n568), 
	.A1N(key_mem[1126]), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U2237 (.Y(n1165), 
	.B1(FE_OFN95_n674), 
	.B0(FE_PHN611_n567), 
	.A1N(FE_PHN1854_key_mem_1127_), 
	.A0N(FE_OFN95_n674));
   OAI2BB2X1 U2238 (.Y(n1160), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN618_n562), 
	.A1N(FE_PHN1777_key_mem_1132_), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U2239 (.Y(n1158), 
	.B1(FE_OFN94_n674), 
	.B0(n560), 
	.A1N(FE_PHN1786_key_mem_1134_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U2240 (.Y(n1156), 
	.B1(FE_OFN94_n674), 
	.B0(n558), 
	.A1N(FE_PHN1810_key_mem_1136_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U2241 (.Y(n1155), 
	.B1(FE_OFN94_n674), 
	.B0(n557), 
	.A1N(FE_PHN1764_key_mem_1137_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U2242 (.Y(n1154), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN614_n556), 
	.A1N(FE_PHN1870_key_mem_1138_), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U2243 (.Y(n1153), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN619_n555), 
	.A1N(key_mem[1139]), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U2244 (.Y(n1152), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN620_n554), 
	.A1N(FE_PHN1819_key_mem_1140_), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U2245 (.Y(n1151), 
	.B1(FE_OFN93_n674), 
	.B0(FE_PHN616_n553), 
	.A1N(FE_PHN1748_key_mem_1141_), 
	.A0N(FE_OFN93_n674));
   OAI2BB2X1 U2246 (.Y(n1150), 
	.B1(FE_OFN94_n674), 
	.B0(n552), 
	.A1N(FE_PHN1846_key_mem_1142_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U2247 (.Y(n1149), 
	.B1(FE_OFN94_n674), 
	.B0(FE_PHN624_n551), 
	.A1N(FE_PHN1874_key_mem_1143_), 
	.A0N(FE_OFN94_n674));
   OAI2BB2X1 U2248 (.Y(n1088), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN389_n618), 
	.A1N(key_mem[1204]), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U2249 (.Y(n1070), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN578_n600), 
	.A1N(FE_PHN1010_key_mem_1222_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U2250 (.Y(n1060), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN421_n590), 
	.A1N(FE_PHN694_key_mem_1232_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U2251 (.Y(n1059), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN419_n589), 
	.A1N(key_mem[1233]), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U2252 (.Y(n1056), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN542_n586), 
	.A1N(FE_PHN968_key_mem_1236_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U2253 (.Y(n1043), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN610_n573), 
	.A1N(FE_PHN779_key_mem_1249_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U2254 (.Y(n1042), 
	.B1(FE_OFN82_n672), 
	.B0(FE_PHN612_n572), 
	.A1N(FE_PHN686_key_mem_1250_), 
	.A0N(FE_OFN82_n672));
   OAI2BB2X1 U2255 (.Y(n1040), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN617_n570), 
	.A1N(FE_PHN688_key_mem_1252_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U2256 (.Y(n1039), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN613_n569), 
	.A1N(FE_PHN1014_key_mem_1253_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U2257 (.Y(n1038), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN605_n568), 
	.A1N(FE_PHN699_key_mem_1254_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U2258 (.Y(n1037), 
	.B1(FE_OFN83_n672), 
	.B0(FE_PHN611_n567), 
	.A1N(FE_PHN1877_key_mem_1255_), 
	.A0N(FE_OFN83_n672));
   OAI2BB2X1 U2259 (.Y(n1032), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN618_n562), 
	.A1N(FE_PHN947_key_mem_1260_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U2260 (.Y(n1030), 
	.B1(FE_OFN81_n672), 
	.B0(n560), 
	.A1N(FE_PHN2831_key_mem_1262_), 
	.A0N(FE_OFN81_n672));
   OAI2BB2X1 U2261 (.Y(n1028), 
	.B1(FE_OFN81_n672), 
	.B0(n558), 
	.A1N(FE_PHN425_key_mem_1264_), 
	.A0N(FE_OFN81_n672));
   OAI2BB2X1 U2262 (.Y(n1027), 
	.B1(n672), 
	.B0(n557), 
	.A1N(FE_PHN700_key_mem_1265_), 
	.A0N(n672));
   OAI2BB2X1 U2263 (.Y(n1026), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN614_n556), 
	.A1N(FE_PHN965_key_mem_1266_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U2264 (.Y(n1025), 
	.B1(n672), 
	.B0(FE_PHN619_n555), 
	.A1N(FE_PHN1780_key_mem_1267_), 
	.A0N(n672));
   OAI2BB2X1 U2265 (.Y(n1024), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN620_n554), 
	.A1N(FE_PHN935_key_mem_1268_), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U2266 (.Y(n1023), 
	.B1(FE_OFN80_n672), 
	.B0(FE_PHN616_n553), 
	.A1N(key_mem[1269]), 
	.A0N(FE_OFN80_n672));
   OAI2BB2X1 U2267 (.Y(n1022), 
	.B1(FE_OFN81_n672), 
	.B0(n552), 
	.A1N(FE_PHN990_key_mem_1270_), 
	.A0N(FE_OFN81_n672));
   OAI2BB2X1 U2268 (.Y(n1021), 
	.B1(FE_OFN81_n672), 
	.B0(FE_PHN624_n551), 
	.A1N(FE_PHN984_key_mem_1271_), 
	.A0N(FE_OFN81_n672));
   OAI2BB2X1 U2269 (.Y(n1344), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN389_n618), 
	.A1N(key_mem[948]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U2270 (.Y(n1326), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN578_n600), 
	.A1N(key_mem[966]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U2271 (.Y(n1316), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN421_n590), 
	.A1N(key_mem[976]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U2272 (.Y(n1315), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN419_n589), 
	.A1N(key_mem[977]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U2273 (.Y(n1312), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN542_n586), 
	.A1N(key_mem[980]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U2274 (.Y(n1299), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN610_n573), 
	.A1N(key_mem[993]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U2275 (.Y(n1298), 
	.B1(FE_OFN77_n676), 
	.B0(FE_PHN612_n572), 
	.A1N(key_mem[994]), 
	.A0N(FE_OFN77_n676));
   OAI2BB2X1 U2276 (.Y(n1296), 
	.B1(n676), 
	.B0(FE_PHN617_n570), 
	.A1N(key_mem[996]), 
	.A0N(n676));
   OAI2BB2X1 U2277 (.Y(n1295), 
	.B1(n676), 
	.B0(FE_PHN613_n569), 
	.A1N(key_mem[997]), 
	.A0N(n676));
   OAI2BB2X1 U2278 (.Y(n1294), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN605_n568), 
	.A1N(key_mem[998]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U2279 (.Y(n1293), 
	.B1(FE_OFN78_n676), 
	.B0(FE_PHN611_n567), 
	.A1N(key_mem[999]), 
	.A0N(FE_OFN78_n676));
   OAI2BB2X1 U2280 (.Y(n1288), 
	.B1(n676), 
	.B0(FE_PHN618_n562), 
	.A1N(key_mem[1004]), 
	.A0N(n676));
   OAI2BB2X1 U2281 (.Y(n1286), 
	.B1(FE_OFN76_n676), 
	.B0(n560), 
	.A1N(key_mem[1006]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U2282 (.Y(n1284), 
	.B1(FE_OFN76_n676), 
	.B0(n558), 
	.A1N(key_mem[1008]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U2283 (.Y(n1283), 
	.B1(FE_OFN76_n676), 
	.B0(n557), 
	.A1N(key_mem[1009]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U2284 (.Y(n1282), 
	.B1(n676), 
	.B0(FE_PHN614_n556), 
	.A1N(key_mem[1010]), 
	.A0N(n676));
   OAI2BB2X1 U2285 (.Y(n1281), 
	.B1(n676), 
	.B0(FE_PHN619_n555), 
	.A1N(key_mem[1011]), 
	.A0N(n676));
   OAI2BB2X1 U2286 (.Y(n1280), 
	.B1(n676), 
	.B0(FE_PHN620_n554), 
	.A1N(key_mem[1012]), 
	.A0N(n676));
   OAI2BB2X1 U2287 (.Y(n1279), 
	.B1(n676), 
	.B0(FE_PHN616_n553), 
	.A1N(key_mem[1013]), 
	.A0N(n676));
   OAI2BB2X1 U2288 (.Y(n1278), 
	.B1(FE_OFN76_n676), 
	.B0(n552), 
	.A1N(key_mem[1014]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U2289 (.Y(n1277), 
	.B1(FE_OFN76_n676), 
	.B0(FE_PHN624_n551), 
	.A1N(key_mem[1015]), 
	.A0N(FE_OFN76_n676));
   OAI2BB2X1 U2290 (.Y(n960), 
	.B1(FE_OFN87_n1), 
	.B0(FE_PHN389_n618), 
	.A1N(key_mem[1332]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U2291 (.Y(n942), 
	.B1(FE_OFN88_n1), 
	.B0(FE_PHN578_n600), 
	.A1N(key_mem[1350]), 
	.A0N(FE_OFN88_n1));
   OAI2BB2X1 U2292 (.Y(n932), 
	.B1(n2624), 
	.B0(FE_PHN421_n590), 
	.A1N(key_mem[1360]), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U2293 (.Y(n931), 
	.B1(n2624), 
	.B0(FE_PHN419_n589), 
	.A1N(key_mem[1361]), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U2294 (.Y(n928), 
	.B1(n2624), 
	.B0(FE_PHN542_n586), 
	.A1N(key_mem[1364]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U2295 (.Y(n915), 
	.B1(n2623), 
	.B0(FE_PHN610_n573), 
	.A1N(key_mem[1377]), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U2296 (.Y(n914), 
	.B1(n2623), 
	.B0(FE_PHN612_n572), 
	.A1N(key_mem[1378]), 
	.A0N(FE_OFN89_n1));
   OAI2BB2X1 U2297 (.Y(n912), 
	.B1(n2623), 
	.B0(FE_PHN617_n570), 
	.A1N(key_mem[1380]), 
	.A0N(n1));
   OAI2BB2X1 U2298 (.Y(n911), 
	.B1(n2623), 
	.B0(FE_PHN613_n569), 
	.A1N(key_mem[1381]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U2299 (.Y(n910), 
	.B1(n2623), 
	.B0(FE_PHN605_n568), 
	.A1N(FE_PHN2836_key_mem_1382_), 
	.A0N(FE_OFN88_n1));
   OAI2BB2X1 U2300 (.Y(n909), 
	.B1(n2622), 
	.B0(FE_PHN611_n567), 
	.A1N(key_mem[1383]), 
	.A0N(FE_OFN86_n1));
   OAI2BB2X1 U2301 (.Y(n904), 
	.B1(n2622), 
	.B0(FE_PHN618_n562), 
	.A1N(key_mem[1388]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U2302 (.Y(n902), 
	.B1(n2622), 
	.B0(n560), 
	.A1N(FE_PHN592_key_mem_1390_), 
	.A0N(FE_OFN85_n1));
   OAI2BB2X1 U2303 (.Y(n900), 
	.B1(n2622), 
	.B0(n558), 
	.A1N(key_mem[1392]), 
	.A0N(FE_OFN85_n1));
   OAI2BB2X1 U2304 (.Y(n899), 
	.B1(n2622), 
	.B0(n557), 
	.A1N(FE_PHN3258_key_mem_1393_), 
	.A0N(n1));
   OAI2BB2X1 U2305 (.Y(n898), 
	.B1(n2622), 
	.B0(FE_PHN614_n556), 
	.A1N(key_mem[1394]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U2306 (.Y(n897), 
	.B1(FE_OFN87_n1), 
	.B0(FE_PHN619_n555), 
	.A1N(key_mem[1395]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U2307 (.Y(n896), 
	.B1(FE_OFN87_n1), 
	.B0(FE_PHN620_n554), 
	.A1N(key_mem[1396]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U2308 (.Y(n895), 
	.B1(FE_OFN87_n1), 
	.B0(FE_PHN616_n553), 
	.A1N(key_mem[1397]), 
	.A0N(FE_OFN87_n1));
   OAI2BB2X1 U2309 (.Y(n894), 
	.B1(FE_OFN85_n1), 
	.B0(n552), 
	.A1N(key_mem[1398]), 
	.A0N(FE_OFN85_n1));
   OAI2BB2X1 U2310 (.Y(n893), 
	.B1(FE_OFN85_n1), 
	.B0(FE_PHN624_n551), 
	.A1N(key_mem[1399]), 
	.A0N(FE_OFN85_n1));
   AOI22X1 U2312 (.Y(n568), 
	.B1(n2649), 
	.B0(key[102]), 
	.A1(n724), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2314 (.Y(n558), 
	.B1(n2644), 
	.B0(key[112]), 
	.A1(n714), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2316 (.Y(n557), 
	.B1(n2644), 
	.B0(key[113]), 
	.A1(n713), 
	.A0(FE_OFN91_n690));
   AOI22X1 U2318 (.Y(n554), 
	.B1(n2642), 
	.B0(key[116]), 
	.A1(n710), 
	.A0(FE_OFN90_n690));
   NOR2BX4 U2319 (.Y(n22), 
	.B(n2877), 
	.AN(round[3]));
   NOR2BX4 U2320 (.Y(n23), 
	.B(n2876), 
	.AN(round[3]));
   INVX1 U2321 (.Y(n2877), 
	.A(round[1]));
   INVX1 U2322 (.Y(n2876), 
	.A(round[0]));
   AOI222X1 U2323 (.Y(n210), 
	.C1(n2806), 
	.C0(key_mem[571]), 
	.B1(n2818), 
	.B0(key_mem[443]), 
	.A1(n2829), 
	.A0(FE_PHN1535_key_mem_699_));
   AOI222X1 U2324 (.Y(n66), 
	.C1(n2800), 
	.C0(key_mem[603]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[475]), 
	.A1(n2823), 
	.A0(FE_PHN1671_key_mem_731_));
   AOI222X1 U2325 (.Y(n350), 
	.C1(n2800), 
	.C0(key_mem[539]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[411]), 
	.A1(n2823), 
	.A0(key_mem[667]));
   AOI222X1 U2326 (.Y(n434), 
	.C1(n2806), 
	.C0(key_mem[635]), 
	.B1(n2818), 
	.B0(key_mem[507]), 
	.A1(n2823), 
	.A0(FE_PHN1552_key_mem_763_));
   AOI222X1 U2327 (.Y(n354), 
	.C1(n2800), 
	.C0(key_mem[538]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[410]), 
	.A1(n2823), 
	.A0(key_mem[666]));
   AOI222X1 U2328 (.Y(n438), 
	.C1(n2806), 
	.C0(key_mem[634]), 
	.B1(n2818), 
	.B0(key_mem[506]), 
	.A1(n2823), 
	.A0(FE_PHN1531_key_mem_762_));
   AOI222X1 U2329 (.Y(n70), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[602]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[474]), 
	.A1(n2823), 
	.A0(FE_PHN1666_key_mem_730_));
   AOI222X1 U2330 (.Y(n214), 
	.C1(n2806), 
	.C0(key_mem[570]), 
	.B1(n2818), 
	.B0(key_mem[442]), 
	.A1(n2829), 
	.A0(FE_PHN1698_key_mem_698_));
   AOI222X1 U2331 (.Y(n218), 
	.C1(n2806), 
	.C0(key_mem[569]), 
	.B1(n2818), 
	.B0(key_mem[441]), 
	.A1(n2829), 
	.A0(FE_PHN1645_key_mem_697_));
   AOI222X1 U2332 (.Y(n358), 
	.C1(n2800), 
	.C0(key_mem[537]), 
	.B1(FE_OFN99_n2811), 
	.B0(FE_PHN3425_key_mem_409_), 
	.A1(n2823), 
	.A0(FE_PHN3214_key_mem_665_));
   AOI222X1 U2333 (.Y(n442), 
	.C1(n2806), 
	.C0(key_mem[633]), 
	.B1(n2818), 
	.B0(key_mem[505]), 
	.A1(n2823), 
	.A0(FE_PHN3196_key_mem_761_));
   AOI222X1 U2334 (.Y(n78), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[601]), 
	.B1(n2817), 
	.B0(key_mem[473]), 
	.A1(n2823), 
	.A0(FE_PHN1528_key_mem_729_));
   AOI222X1 U2335 (.Y(n82), 
	.C1(n2800), 
	.C0(key_mem[600]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[472]), 
	.A1(n2823), 
	.A0(FE_PHN1642_key_mem_728_));
   AOI222X1 U2336 (.Y(n362), 
	.C1(n2800), 
	.C0(key_mem[536]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[408]), 
	.A1(n2823), 
	.A0(FE_PHN1512_key_mem_664_));
   AOI222X1 U2337 (.Y(n446), 
	.C1(n2800), 
	.C0(key_mem[632]), 
	.B1(FE_OFN99_n2811), 
	.B0(FE_PHN2826_key_mem_504_), 
	.A1(n2824), 
	.A0(FE_PHN772_key_mem_760_));
   AOI222X1 U2338 (.Y(n418), 
	.C1(n2806), 
	.C0(key_mem[639]), 
	.B1(n2818), 
	.B0(FE_PHN3221_key_mem_511_), 
	.A1(n2823), 
	.A0(FE_PHN762_key_mem_767_));
   AOI222X1 U2339 (.Y(n422), 
	.C1(n2806), 
	.C0(key_mem[638]), 
	.B1(n2818), 
	.B0(key_mem[510]), 
	.A1(n2823), 
	.A0(FE_PHN756_key_mem_766_));
   AOI222X1 U2340 (.Y(n426), 
	.C1(n2806), 
	.C0(key_mem[637]), 
	.B1(n2818), 
	.B0(key_mem[509]), 
	.A1(n2823), 
	.A0(FE_PHN1602_key_mem_765_));
   AOI222X1 U2341 (.Y(n62), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[604]), 
	.B1(n2817), 
	.B0(key_mem[476]), 
	.A1(n2823), 
	.A0(FE_PHN1746_key_mem_732_));
   AOI222X1 U2342 (.Y(n222), 
	.C1(n2806), 
	.C0(key_mem[568]), 
	.B1(n2818), 
	.B0(key_mem[440]), 
	.A1(n2829), 
	.A0(FE_PHN1771_key_mem_696_));
   AOI222X1 U2343 (.Y(n190), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[575]), 
	.B1(n2818), 
	.B0(key_mem[447]), 
	.A1(n2828), 
	.A0(FE_PHN758_key_mem_703_));
   AOI222X1 U2344 (.Y(n194), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[574]), 
	.B1(n2818), 
	.B0(key_mem[446]), 
	.A1(n2828), 
	.A0(FE_PHN1516_key_mem_702_));
   AOI222X1 U2345 (.Y(n198), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[573]), 
	.B1(n2818), 
	.B0(key_mem[445]), 
	.A1(n2828), 
	.A0(FE_PHN1656_key_mem_701_));
   AOI222X1 U2346 (.Y(n202), 
	.C1(n2800), 
	.C0(key_mem[572]), 
	.B1(n2818), 
	.B0(key_mem[444]), 
	.A1(n2828), 
	.A0(FE_PHN1483_key_mem_700_));
   AOI222X1 U2347 (.Y(n346), 
	.C1(n2800), 
	.C0(key_mem[540]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[412]), 
	.A1(n2827), 
	.A0(key_mem[668]));
   AOI222X1 U2348 (.Y(n430), 
	.C1(n2806), 
	.C0(key_mem[636]), 
	.B1(n2818), 
	.B0(key_mem[508]), 
	.A1(n2823), 
	.A0(FE_PHN1765_key_mem_764_));
   AOI222X1 U2349 (.Y(n330), 
	.C1(n2800), 
	.C0(FE_PHN3410_key_mem_543_), 
	.B1(FE_OFN99_n2811), 
	.B0(FE_PHN3184_key_mem_415_), 
	.A1(n2827), 
	.A0(FE_PHN1706_key_mem_671_));
   AOI222X1 U2350 (.Y(n334), 
	.C1(n2800), 
	.C0(key_mem[542]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[414]), 
	.A1(n2827), 
	.A0(FE_PHN1569_key_mem_670_));
   AOI222X1 U2351 (.Y(n342), 
	.C1(n2800), 
	.C0(key_mem[541]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[413]), 
	.A1(n2827), 
	.A0(key_mem[669]));
   AOI222X1 U2352 (.Y(n38), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[610]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[482]), 
	.A1(n2823), 
	.A0(FE_PHN1824_key_mem_738_));
   AOI222X1 U2353 (.Y(n34), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[611]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[483]), 
	.A1(n2823), 
	.A0(FE_PHN1692_key_mem_739_));
   AOI222X1 U2354 (.Y(n19), 
	.C1(n2800), 
	.C0(key_mem[521]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[393]), 
	.A1(n2823), 
	.A0(FE_PHN1481_key_mem_649_));
   AOI222X1 U2355 (.Y(n42), 
	.C1(n2800), 
	.C0(key_mem[609]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[481]), 
	.A1(n2823), 
	.A0(FE_PHN1804_key_mem_737_));
   AOI222X1 U2356 (.Y(n46), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[608]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[480]), 
	.A1(n2823), 
	.A0(FE_PHN1520_key_mem_736_));
   AOI222X1 U2357 (.Y(n54), 
	.C1(n2800), 
	.C0(key_mem[606]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[478]), 
	.A1(n2823), 
	.A0(FE_PHN1680_key_mem_734_));
   AOI222X1 U2358 (.Y(n58), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[605]), 
	.B1(n2817), 
	.B0(key_mem[477]), 
	.A1(n2823), 
	.A0(FE_PHN1587_key_mem_733_));
   AOI222X1 U2359 (.Y(n50), 
	.C1(n2800), 
	.C0(key_mem[607]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[479]), 
	.A1(n2823), 
	.A0(FE_PHN1596_key_mem_735_));
   AOI222X1 U2360 (.Y(n493), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[906]), 
	.B1(n2775), 
	.B0(key_mem[778]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN3303_key_mem_1034_));
   AOI222X1 U2361 (.Y(n337), 
	.C1(FE_OFN105_n2763), 
	.C0(FE_PHN3434_key_mem_898_), 
	.B1(n2780), 
	.B0(FE_PHN3412_key_mem_770_), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN3239_key_mem_1026_));
   AOI222X1 U2362 (.Y(n321), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[929]), 
	.B1(n2780), 
	.B0(key_mem[801]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1832_key_mem_1057_));
   AOI222X1 U2363 (.Y(n293), 
	.C1(n2769), 
	.C0(key_mem[899]), 
	.B1(n2781), 
	.B0(key_mem[771]), 
	.A1(FE_OFN104_n27), 
	.A0(key_mem[1027]));
   AOI222X1 U2364 (.Y(n317), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[930]), 
	.B1(n2780), 
	.B0(key_mem[802]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1743_key_mem_1058_));
   AOI222X1 U2365 (.Y(n469), 
	.C1(n2769), 
	.C0(key_mem[1011]), 
	.B1(n2775), 
	.B0(key_mem[883]), 
	.A1(FE_OFN103_n27), 
	.A0(key_mem[1139]));
   AOI222X1 U2366 (.Y(n389), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[914]), 
	.B1(n2775), 
	.B0(key_mem[786]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1719_key_mem_1042_));
   AOI222X1 U2367 (.Y(n473), 
	.C1(n2769), 
	.C0(key_mem[1010]), 
	.B1(n2775), 
	.B0(key_mem[882]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1870_key_mem_1138_));
   AOI222X1 U2368 (.Y(n105), 
	.C1(n2773), 
	.C0(key_mem[978]), 
	.B1(n2775), 
	.B0(key_mem[850]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1871_key_mem_1106_));
   AOI222X1 U2369 (.Y(n245), 
	.C1(n2770), 
	.C0(key_mem[946]), 
	.B1(n2781), 
	.B0(key_mem[818]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1773_key_mem_1074_));
   AOI222X1 U2370 (.Y(n393), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[913]), 
	.B1(n2775), 
	.B0(key_mem[785]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1840_key_mem_1041_));
   AOI222X1 U2371 (.Y(n145), 
	.C1(FE_OFN105_n2763), 
	.C0(FE_PHN3433_key_mem_969_), 
	.B1(n2784), 
	.B0(FE_PHN3186_key_mem_841_), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1799_key_mem_1097_));
   AOI222X1 U2372 (.Y(n513), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[1001]), 
	.B1(n2775), 
	.B0(key_mem[873]), 
	.A1(FE_OFN103_n27), 
	.A0(key_mem[1129]));
   AOI222X1 U2373 (.Y(n477), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[1009]), 
	.B1(n2775), 
	.B0(key_mem[881]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1764_key_mem_1137_));
   AOI222X1 U2374 (.Y(n109), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[977]), 
	.B1(n2784), 
	.B0(key_mem[849]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1745_key_mem_1105_));
   AOI222X1 U2375 (.Y(n253), 
	.C1(n2769), 
	.C0(key_mem[945]), 
	.B1(n2781), 
	.B0(key_mem[817]), 
	.A1(FE_OFN104_n27), 
	.A0(key_mem[1073]));
   AOI222X1 U2376 (.Y(n113), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[976]), 
	.B1(n2784), 
	.B0(key_mem[848]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1821_key_mem_1104_));
   AOI222X1 U2377 (.Y(n73), 
	.C1(n2773), 
	.C0(key_mem[904]), 
	.B1(n2775), 
	.B0(key_mem[776]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1713_key_mem_1032_));
   AOI222X1 U2378 (.Y(n257), 
	.C1(n2769), 
	.C0(key_mem[944]), 
	.B1(n2781), 
	.B0(key_mem[816]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1861_key_mem_1072_));
   AOI222X1 U2379 (.Y(n397), 
	.C1(n2766), 
	.C0(key_mem[912]), 
	.B1(n2775), 
	.B0(key_mem[784]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1881_key_mem_1040_));
   AOI222X1 U2380 (.Y(n481), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[1008]), 
	.B1(n2775), 
	.B0(key_mem[880]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1810_key_mem_1136_));
   AOI222X1 U2381 (.Y(n289), 
	.C1(n2769), 
	.C0(key_mem[936]), 
	.B1(n2781), 
	.B0(key_mem[808]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1852_key_mem_1064_));
   AOI222X1 U2382 (.Y(n517), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[1000]), 
	.B1(n2775), 
	.B0(key_mem[872]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1816_key_mem_1128_));
   AOI222X1 U2383 (.Y(n365), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[919]), 
	.B1(n2775), 
	.B0(FE_PHN3198_key_mem_791_), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1761_key_mem_1047_));
   AOI222X1 U2384 (.Y(n453), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[1015]), 
	.B1(n2775), 
	.B0(key_mem[887]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1874_key_mem_1143_));
   AOI222X1 U2385 (.Y(n85), 
	.C1(n2773), 
	.C0(key_mem[983]), 
	.B1(n2775), 
	.B0(key_mem[855]), 
	.A1(FE_OFN103_n27), 
	.A0(key_mem[1111]));
   AOI222X1 U2386 (.Y(n225), 
	.C1(n2770), 
	.C0(key_mem[951]), 
	.B1(n2781), 
	.B0(key_mem[823]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1829_key_mem_1079_));
   AOI222X1 U2387 (.Y(n153), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[967]), 
	.B1(n2784), 
	.B0(key_mem[839]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1778_key_mem_1095_));
   AOI222X1 U2388 (.Y(n89), 
	.C1(n2773), 
	.C0(key_mem[982]), 
	.B1(n2775), 
	.B0(key_mem[854]), 
	.A1(FE_OFN104_n27), 
	.A0(key_mem[1110]));
   AOI222X1 U2389 (.Y(n229), 
	.C1(n2770), 
	.C0(key_mem[950]), 
	.B1(n2781), 
	.B0(key_mem[822]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1866_key_mem_1078_));
   AOI222X1 U2390 (.Y(n369), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[918]), 
	.B1(n2775), 
	.B0(key_mem[790]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1905_key_mem_1046_));
   AOI222X1 U2391 (.Y(n457), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[1014]), 
	.B1(n2775), 
	.B0(key_mem[886]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1846_key_mem_1142_));
   AOI222X1 U2392 (.Y(n93), 
	.C1(n2773), 
	.C0(key_mem[981]), 
	.B1(n2775), 
	.B0(key_mem[853]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1787_key_mem_1109_));
   AOI222X1 U2393 (.Y(n233), 
	.C1(n2770), 
	.C0(key_mem[949]), 
	.B1(n2781), 
	.B0(key_mem[821]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1789_key_mem_1077_));
   AOI222X1 U2394 (.Y(n373), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[917]), 
	.B1(n2775), 
	.B0(key_mem[789]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1880_key_mem_1045_));
   AOI222X1 U2395 (.Y(n129), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[973]), 
	.B1(n2784), 
	.B0(key_mem[845]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1893_key_mem_1101_));
   AOI222X1 U2396 (.Y(n237), 
	.C1(n2770), 
	.C0(key_mem[948]), 
	.B1(n2781), 
	.B0(key_mem[820]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1798_key_mem_1076_));
   AOI222X1 U2397 (.Y(n385), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[915]), 
	.B1(n2775), 
	.B0(key_mem[787]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1833_key_mem_1043_));
   AOI222X1 U2398 (.Y(n137), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[971]), 
	.B1(n2784), 
	.B0(key_mem[843]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1859_key_mem_1099_));
   AOI222X1 U2399 (.Y(n381), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[897]), 
	.B1(n2775), 
	.B0(key_mem[769]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1882_key_mem_1025_));
   AOI222X1 U2400 (.Y(n325), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[928]), 
	.B1(n2780), 
	.B0(key_mem[800]), 
	.A1(FE_OFN104_n27), 
	.A0(key_mem[1056]));
   AOI222X1 U2401 (.Y(n377), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[916]), 
	.B1(n2775), 
	.B0(key_mem[788]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1894_key_mem_1044_));
   AOI222X1 U2402 (.Y(n465), 
	.C1(n2769), 
	.C0(key_mem[1012]), 
	.B1(n2775), 
	.B0(key_mem[884]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1819_key_mem_1140_));
   AOI222X1 U2403 (.Y(n101), 
	.C1(n2773), 
	.C0(key_mem[979]), 
	.B1(n2775), 
	.B0(key_mem[851]), 
	.A1(FE_OFN103_n27), 
	.A0(key_mem[1107]));
   AOI222X1 U2404 (.Y(n117), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[903]), 
	.B1(n2784), 
	.B0(key_mem[775]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1760_key_mem_1031_));
   AOI222X1 U2405 (.Y(n121), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[975]), 
	.B1(n2784), 
	.B0(key_mem[847]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1855_key_mem_1103_));
   AOI222X1 U2406 (.Y(n405), 
	.C1(n2766), 
	.C0(key_mem[910]), 
	.B1(n2775), 
	.B0(key_mem[782]), 
	.A1(FE_OFN103_n27), 
	.A0(key_mem[1038]));
   AOI222X1 U2407 (.Y(n461), 
	.C1(n2769), 
	.C0(key_mem[1013]), 
	.B1(n2775), 
	.B0(key_mem[885]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1748_key_mem_1141_));
   AOI222X1 U2408 (.Y(n273), 
	.C1(n2769), 
	.C0(key_mem[940]), 
	.B1(n2781), 
	.B0(key_mem[812]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1891_key_mem_1068_));
   AOI222X1 U2409 (.Y(n173), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[963]), 
	.B1(n2781), 
	.B0(FE_PHN1469_key_mem_835_), 
	.A1(FE_OFN104_n27), 
	.A0(key_mem[1091]));
   AOI222X1 U2410 (.Y(n449), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[907]), 
	.B1(n2775), 
	.B0(key_mem[779]), 
	.A1(FE_OFN103_n27), 
	.A0(key_mem[1035]));
   AOI222X1 U2411 (.Y(n141), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[970]), 
	.B1(n2784), 
	.B0(key_mem[842]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1756_key_mem_1098_));
   AOI222X1 U2412 (.Y(n149), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[968]), 
	.B1(n2784), 
	.B0(FE_PHN1491_key_mem_840_), 
	.A1(FE_OFN104_n27), 
	.A0(key_mem[1096]));
   AOI222X1 U2413 (.Y(n401), 
	.C1(n2766), 
	.C0(key_mem[911]), 
	.B1(n2775), 
	.B0(FE_PHN3234_key_mem_783_), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1888_key_mem_1039_));
   AOI222X1 U2414 (.Y(n125), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[974]), 
	.B1(n2784), 
	.B0(FE_PHN2789_key_mem_846_), 
	.A1(FE_OFN104_n27), 
	.A0(key_mem[1102]));
   AOI222X1 U2415 (.Y(n409), 
	.C1(n2766), 
	.C0(key_mem[909]), 
	.B1(n2775), 
	.B0(key_mem[781]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1788_key_mem_1037_));
   AOI222X1 U2416 (.Y(n133), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[972]), 
	.B1(n2784), 
	.B0(key_mem[844]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1887_key_mem_1100_));
   AOI222X1 U2417 (.Y(n533), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[996]), 
	.B1(n2775), 
	.B0(key_mem[868]), 
	.A1(FE_OFN103_n27), 
	.A0(key_mem[1124]));
   AOI222X1 U2418 (.Y(n97), 
	.C1(n2773), 
	.C0(key_mem[980]), 
	.B1(n2775), 
	.B0(key_mem[852]), 
	.A1(FE_OFN103_n27), 
	.A0(key_mem[1108]));
   AOI222X1 U2419 (.Y(n241), 
	.C1(n2770), 
	.C0(key_mem[947]), 
	.B1(n2781), 
	.B0(key_mem[819]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1712_key_mem_1075_));
   AOI222X1 U2420 (.Y(n509), 
	.C1(FE_OFN105_n2763), 
	.C0(FE_PHN3426_key_mem_1002_), 
	.B1(n2775), 
	.B0(FE_PHN3421_key_mem_874_), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN3307_key_mem_1130_));
   AOI222X1 U2421 (.Y(n285), 
	.C1(n2769), 
	.C0(key_mem[937]), 
	.B1(n2781), 
	.B0(key_mem[809]), 
	.A1(FE_OFN104_n27), 
	.A0(key_mem[1065]));
   AOI222X1 U2422 (.Y(n185), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[960]), 
	.B1(n2781), 
	.B0(key_mem[832]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1869_key_mem_1088_));
   AOI222X1 U2423 (.Y(n521), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[999]), 
	.B1(n2775), 
	.B0(key_mem[871]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1854_key_mem_1127_));
   AOI222X1 U2424 (.Y(n261), 
	.C1(n2769), 
	.C0(key_mem[943]), 
	.B1(n2781), 
	.B0(key_mem[815]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1889_key_mem_1071_));
   AOI222X1 U2425 (.Y(n157), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[966]), 
	.B1(n2781), 
	.B0(key_mem[838]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1863_key_mem_1094_));
   AOI222X1 U2426 (.Y(n525), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[998]), 
	.B1(n2775), 
	.B0(key_mem[870]), 
	.A1(FE_OFN104_n27), 
	.A0(key_mem[1126]));
   AOI222X1 U2427 (.Y(n265), 
	.C1(n2769), 
	.C0(key_mem[942]), 
	.B1(n2781), 
	.B0(key_mem[814]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1758_key_mem_1070_));
   AOI222X1 U2428 (.Y(n165), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[965]), 
	.B1(n2781), 
	.B0(key_mem[837]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1790_key_mem_1093_));
   AOI222X1 U2429 (.Y(n529), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[997]), 
	.B1(n2775), 
	.B0(key_mem[869]), 
	.A1(FE_OFN103_n27), 
	.A0(key_mem[1125]));
   AOI222X1 U2430 (.Y(n269), 
	.C1(n2769), 
	.C0(key_mem[941]), 
	.B1(n2781), 
	.B0(key_mem[813]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1867_key_mem_1069_));
   AOI222X1 U2431 (.Y(n169), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[964]), 
	.B1(n2781), 
	.B0(key_mem[836]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1841_key_mem_1092_));
   AOI222X1 U2432 (.Y(n413), 
	.C1(n2766), 
	.C0(key_mem[908]), 
	.B1(n2775), 
	.B0(key_mem[780]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1811_key_mem_1036_));
   AOI222X1 U2433 (.Y(n309), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[932]), 
	.B1(n2780), 
	.B0(key_mem[804]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1872_key_mem_1060_));
   AOI222X1 U2434 (.Y(n501), 
	.C1(n2769), 
	.C0(key_mem[1004]), 
	.B1(n2775), 
	.B0(key_mem[876]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1777_key_mem_1132_));
   AOI222X1 U2435 (.Y(n277), 
	.C1(n2769), 
	.C0(key_mem[939]), 
	.B1(n2781), 
	.B0(FE_PHN1560_key_mem_811_), 
	.A1(FE_OFN104_n27), 
	.A0(key_mem[1067]));
   AOI222X1 U2436 (.Y(n177), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[962]), 
	.B1(n2781), 
	.B0(key_mem[834]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1830_key_mem_1090_));
   AOI222X1 U2437 (.Y(n537), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[896]), 
	.B1(n2775), 
	.B0(key_mem[768]), 
	.A1(FE_OFN104_n27), 
	.A0(key_mem[1024]));
   AOI222X1 U2438 (.Y(n297), 
	.C1(n2769), 
	.C0(key_mem[935]), 
	.B1(n2781), 
	.B0(key_mem[807]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN954_key_mem_1063_));
   AOI222X1 U2439 (.Y(n485), 
	.C1(FE_OFN105_n2763), 
	.C0(FE_PHN3431_key_mem_1007_), 
	.B1(n2775), 
	.B0(FE_PHN3236_key_mem_879_), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1791_key_mem_1135_));
   AOI222X1 U2440 (.Y(n161), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[902]), 
	.B1(n2781), 
	.B0(key_mem[774]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1862_key_mem_1030_));
   AOI222X1 U2441 (.Y(n301), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[934]), 
	.B1(n2780), 
	.B0(FE_PHN1532_key_mem_806_), 
	.A1(FE_OFN104_n27), 
	.A0(key_mem[1062]));
   AOI222X1 U2442 (.Y(n489), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[1006]), 
	.B1(n2775), 
	.B0(key_mem[878]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1786_key_mem_1134_));
   AOI222X1 U2443 (.Y(n205), 
	.C1(n2770), 
	.C0(key_mem[901]), 
	.B1(n2781), 
	.B0(key_mem[773]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1892_key_mem_1029_));
   AOI222X1 U2444 (.Y(n305), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[933]), 
	.B1(n2780), 
	.B0(key_mem[805]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1873_key_mem_1061_));
   AOI222X1 U2445 (.Y(n497), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[1005]), 
	.B1(n2775), 
	.B0(key_mem[877]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1822_key_mem_1133_));
   AOI222X1 U2446 (.Y(n249), 
	.C1(n2770), 
	.C0(key_mem[900]), 
	.B1(n2781), 
	.B0(key_mem[772]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1853_key_mem_1028_));
   AOI222X1 U2447 (.Y(n313), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[931]), 
	.B1(n2780), 
	.B0(key_mem[803]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1839_key_mem_1059_));
   AOI222X1 U2448 (.Y(n505), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[1003]), 
	.B1(n2775), 
	.B0(key_mem[875]), 
	.A1(FE_OFN103_n27), 
	.A0(key_mem[1131]));
   AOI222X1 U2449 (.Y(n281), 
	.C1(n2769), 
	.C0(key_mem[938]), 
	.B1(n2781), 
	.B0(key_mem[810]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1813_key_mem_1066_));
   AOI222X1 U2450 (.Y(n181), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[961]), 
	.B1(n2781), 
	.B0(key_mem[833]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1701_key_mem_1089_));
   NAND4X1 U2451 (.Y(round_key[98]), 
	.D(n39), 
	.C(n38), 
	.B(n37), 
	.A(n36));
   AOI22X1 U2452 (.Y(n36), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1378]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN686_key_mem_1250_));
   AOI222X1 U2453 (.Y(n39), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[226]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[98]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1659_key_mem_354_));
   AOI222X1 U2454 (.Y(n37), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[994]), 
	.B1(n2775), 
	.B0(key_mem[866]), 
	.A1(FE_OFN104_n27), 
	.A0(key_mem[1122]));
   NAND4X1 U2455 (.Y(round_key[9]), 
	.D(n20), 
	.C(n19), 
	.B(n18), 
	.A(n17));
   AOI22X1 U2456 (.Y(n17), 
	.B1(FE_OFN102_n31), 
	.B0(FE_PHN3205_key_mem_1289_), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN587_key_mem_1161_));
   AOI222X1 U2457 (.Y(n20), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[137]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[9]), 
	.A1(n21), 
	.A0(FE_PHN1688_key_mem_265_));
   AOI222X1 U2458 (.Y(n18), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[905]), 
	.B1(n2775), 
	.B0(FE_PHN3417_key_mem_777_), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN2838_key_mem_1033_));
   NAND4X1 U2459 (.Y(round_key[97]), 
	.D(n43), 
	.C(n42), 
	.B(n41), 
	.A(n40));
   AOI22X1 U2460 (.Y(n40), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1377]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN779_key_mem_1249_));
   AOI222X1 U2461 (.Y(n43), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[225]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[97]), 
	.A1(n21), 
	.A0(FE_PHN1793_key_mem_353_));
   AOI222X1 U2462 (.Y(n41), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[993]), 
	.B1(n2775), 
	.B0(key_mem[865]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1850_key_mem_1121_));
   NAND4X1 U2463 (.Y(n690), 
	.D(n2874), 
	.C(n2873), 
	.B(n2872), 
	.A(FE_PHN411_n6));
   INVX1 U2464 (.Y(n2878), 
	.A(round[2]));
   AND3X4 U2465 (.Y(n21), 
	.C(round[3]), 
	.B(n2877), 
	.A(n2876));
   NOR3X1 U2466 (.Y(n540), 
	.C(round[1]), 
	.B(round[3]), 
	.A(round[2]));
   NAND4X1 U2467 (.Y(round_key[10]), 
	.D(n495), 
	.C(n494), 
	.B(n493), 
	.A(n492));
   AOI22X1 U2468 (.Y(n492), 
	.B1(n31), 
	.B0(FE_PHN3285_key_mem_1290_), 
	.A1(n30), 
	.A0(FE_PHN429_key_mem_1162_));
   AOI222X1 U2469 (.Y(n495), 
	.C1(n23), 
	.C0(FE_PHN3428_key_mem_138_), 
	.B1(n22), 
	.B0(FE_PHN3206_key_mem_10_), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1697_key_mem_266_));
   AOI222X1 U2470 (.Y(n494), 
	.C1(n2800), 
	.C0(FE_PHN3416_key_mem_522_), 
	.B1(FE_OFN99_n2811), 
	.B0(FE_PHN3430_key_mem_394_), 
	.A1(n2823), 
	.A0(FE_PHN2832_key_mem_650_));
   NAND4X1 U2471 (.Y(round_key[2]), 
	.D(n339), 
	.C(n338), 
	.B(n337), 
	.A(n336));
   AOI22X1 U2472 (.Y(n336), 
	.B1(n31), 
	.B0(FE_PHN2825_key_mem_1282_), 
	.A1(n30), 
	.A0(FE_PHN357_key_mem_1154_));
   AOI222X1 U2473 (.Y(n339), 
	.C1(n23), 
	.C0(FE_PHN3429_key_mem_130_), 
	.B1(n22), 
	.B0(FE_PHN3248_key_mem_2_), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1703_key_mem_258_));
   AOI222X1 U2474 (.Y(n338), 
	.C1(n2800), 
	.C0(FE_PHN3437_key_mem_514_), 
	.B1(FE_OFN99_n2811), 
	.B0(FE_PHN3226_key_mem_386_), 
	.A1(n2827), 
	.A0(FE_PHN1502_key_mem_642_));
   NAND4X1 U2475 (.Y(round_key[33]), 
	.D(n323), 
	.C(n322), 
	.B(n321), 
	.A(n320));
   AOI22X1 U2476 (.Y(n320), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1313]), 
	.A1(FE_OFN101_n30), 
	.A0(key_mem[1185]));
   AOI222X1 U2477 (.Y(n323), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[161]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[33]), 
	.A1(n21), 
	.A0(FE_PHN1492_key_mem_289_));
   AOI222X1 U2478 (.Y(n322), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[545]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[417]), 
	.A1(n2827), 
	.A0(FE_PHN1694_key_mem_673_));
   NAND4X1 U2479 (.Y(round_key[3]), 
	.D(n295), 
	.C(n294), 
	.B(n293), 
	.A(n292));
   AOI22X1 U2480 (.Y(n292), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1283]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN1023_key_mem_1155_));
   AOI222X1 U2481 (.Y(n295), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[131]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[3]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1546_key_mem_259_));
   AOI222X1 U2482 (.Y(n294), 
	.C1(n2806), 
	.C0(key_mem[515]), 
	.B1(n2817), 
	.B0(key_mem[387]), 
	.A1(n2828), 
	.A0(FE_PHN1615_key_mem_643_));
   NAND4X1 U2483 (.Y(round_key[34]), 
	.D(n319), 
	.C(n318), 
	.B(n317), 
	.A(n316));
   AOI22X1 U2484 (.Y(n316), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1314]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN1015_key_mem_1186_));
   AOI222X1 U2485 (.Y(n319), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[162]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[34]), 
	.A1(n21), 
	.A0(FE_PHN1573_key_mem_290_));
   AOI222X1 U2486 (.Y(n318), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[546]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[418]), 
	.A1(n2827), 
	.A0(FE_PHN1641_key_mem_674_));
   NAND4X1 U2487 (.Y(round_key[115]), 
	.D(n471), 
	.C(n470), 
	.B(n469), 
	.A(n468));
   AOI22X1 U2488 (.Y(n468), 
	.B1(n31), 
	.B0(key_mem[1395]), 
	.A1(n30), 
	.A0(FE_PHN1780_key_mem_1267_));
   AOI222X1 U2489 (.Y(n471), 
	.C1(n23), 
	.C0(key_mem[243]), 
	.B1(n22), 
	.B0(key_mem[115]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN915_key_mem_371_));
   AOI222X1 U2490 (.Y(n470), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[627]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[499]), 
	.A1(n2824), 
	.A0(FE_PHN1828_key_mem_755_));
   NAND4X1 U2491 (.Y(round_key[18]), 
	.D(n391), 
	.C(n390), 
	.B(n389), 
	.A(n388));
   AOI22X1 U2492 (.Y(n388), 
	.B1(n31), 
	.B0(FE_PHN2823_key_mem_1298_), 
	.A1(n30), 
	.A0(FE_PHN582_key_mem_1170_));
   AOI222X1 U2493 (.Y(n391), 
	.C1(n23), 
	.C0(key_mem[146]), 
	.B1(n22), 
	.B0(FE_PHN3194_key_mem_18_), 
	.A1(n21), 
	.A0(FE_PHN1639_key_mem_274_));
   AOI222X1 U2494 (.Y(n390), 
	.C1(n2800), 
	.C0(key_mem[530]), 
	.B1(FE_OFN99_n2811), 
	.B0(FE_PHN3195_key_mem_402_), 
	.A1(n2823), 
	.A0(FE_PHN1505_key_mem_658_));
   NAND4X1 U2495 (.Y(round_key[114]), 
	.D(n475), 
	.C(n474), 
	.B(n473), 
	.A(n472));
   AOI22X1 U2496 (.Y(n472), 
	.B1(n31), 
	.B0(key_mem[1394]), 
	.A1(n30), 
	.A0(FE_PHN965_key_mem_1266_));
   AOI222X1 U2497 (.Y(n475), 
	.C1(n23), 
	.C0(key_mem[242]), 
	.B1(n22), 
	.B0(key_mem[114]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1644_key_mem_370_));
   AOI222X1 U2498 (.Y(n474), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[626]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[498]), 
	.A1(n2824), 
	.A0(FE_PHN1536_key_mem_754_));
   NAND4X1 U2499 (.Y(round_key[82]), 
	.D(n107), 
	.C(n106), 
	.B(n105), 
	.A(n104));
   AOI22X1 U2500 (.Y(n104), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1362]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN777_key_mem_1234_));
   AOI222X1 U2501 (.Y(n107), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[210]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[82]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1637_key_mem_338_));
   AOI222X1 U2502 (.Y(n106), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[594]), 
	.B1(n2817), 
	.B0(key_mem[466]), 
	.A1(n2823), 
	.A0(FE_PHN1519_key_mem_722_));
   NAND4X1 U2503 (.Y(round_key[50]), 
	.D(n247), 
	.C(n246), 
	.B(n245), 
	.A(n244));
   AOI22X1 U2504 (.Y(n244), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1330]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN992_key_mem_1202_));
   AOI222X1 U2505 (.Y(n247), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[178]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[50]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1559_key_mem_306_));
   AOI222X1 U2506 (.Y(n246), 
	.C1(n2806), 
	.C0(key_mem[562]), 
	.B1(n2818), 
	.B0(key_mem[434]), 
	.A1(n2829), 
	.A0(FE_PHN1506_key_mem_690_));
   NAND4X1 U2507 (.Y(round_key[17]), 
	.D(n395), 
	.C(n394), 
	.B(n393), 
	.A(n392));
   AOI22X1 U2508 (.Y(n392), 
	.B1(n31), 
	.B0(FE_PHN2837_key_mem_1297_), 
	.A1(n30), 
	.A0(FE_PHN1792_key_mem_1169_));
   AOI222X1 U2509 (.Y(n395), 
	.C1(n23), 
	.C0(key_mem[145]), 
	.B1(n22), 
	.B0(key_mem[17]), 
	.A1(n21), 
	.A0(FE_PHN1542_key_mem_273_));
   AOI222X1 U2510 (.Y(n394), 
	.C1(n2800), 
	.C0(key_mem[529]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[401]), 
	.A1(n2823), 
	.A0(FE_PHN754_key_mem_657_));
   NAND4X1 U2511 (.Y(round_key[73]), 
	.D(n147), 
	.C(n146), 
	.B(n145), 
	.A(n144));
   AOI22X1 U2512 (.Y(n144), 
	.B1(FE_OFN102_n31), 
	.B0(FE_PHN2841_key_mem_1353_), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN594_key_mem_1225_));
   AOI222X1 U2513 (.Y(n147), 
	.C1(FE_OFN109_n23), 
	.C0(FE_PHN3424_key_mem_201_), 
	.B1(FE_OFN106_n22), 
	.B0(FE_PHN3189_key_mem_73_), 
	.A1(n21), 
	.A0(FE_PHN1627_key_mem_329_));
   AOI222X1 U2514 (.Y(n146), 
	.C1(FE_OFN100_n2800), 
	.C0(FE_PHN3414_key_mem_585_), 
	.B1(FE_OFN99_n2811), 
	.B0(FE_PHN3197_key_mem_457_), 
	.A1(n2823), 
	.A0(FE_PHN1820_key_mem_713_));
   NAND4X1 U2516 (.Y(round_key[105]), 
	.D(n515), 
	.C(n514), 
	.B(n513), 
	.A(n512));
   AOI22X1 U2517 (.Y(n512), 
	.B1(n31), 
	.B0(key_mem[1385]), 
	.A1(n30), 
	.A0(FE_PHN583_key_mem_1257_));
   AOI222X1 U2518 (.Y(n515), 
	.C1(n23), 
	.C0(key_mem[233]), 
	.B1(n22), 
	.B0(key_mem[105]), 
	.A1(n21), 
	.A0(FE_PHN1595_key_mem_361_));
   AOI222X1 U2519 (.Y(n514), 
	.C1(n2800), 
	.C0(key_mem[617]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[489]), 
	.A1(n2823), 
	.A0(key_mem[745]));
   NAND4X1 U2520 (.Y(round_key[113]), 
	.D(n479), 
	.C(n478), 
	.B(n477), 
	.A(n476));
   AOI22X1 U2521 (.Y(n476), 
	.B1(n31), 
	.B0(FE_PHN3258_key_mem_1393_), 
	.A1(n30), 
	.A0(FE_PHN700_key_mem_1265_));
   AOI222X1 U2522 (.Y(n479), 
	.C1(n23), 
	.C0(key_mem[241]), 
	.B1(n22), 
	.B0(key_mem[113]), 
	.A1(n21), 
	.A0(FE_PHN1605_key_mem_369_));
   AOI222X1 U2523 (.Y(n478), 
	.C1(n2800), 
	.C0(key_mem[625]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[497]), 
	.A1(n2824), 
	.A0(FE_PHN2824_key_mem_753_));
   NAND4X1 U2524 (.Y(round_key[81]), 
	.D(n111), 
	.C(n110), 
	.B(n109), 
	.A(n108));
   AOI22X1 U2525 (.Y(n108), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1361]), 
	.A1(FE_OFN101_n30), 
	.A0(key_mem[1233]));
   AOI222X1 U2526 (.Y(n111), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[209]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[81]), 
	.A1(n21), 
	.A0(FE_PHN1533_key_mem_337_));
   AOI222X1 U2527 (.Y(n110), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[593]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[465]), 
	.A1(n2823), 
	.A0(FE_PHN1718_key_mem_721_));
   NAND4X1 U2528 (.Y(round_key[49]), 
	.D(n255), 
	.C(n254), 
	.B(n253), 
	.A(n252));
   AOI22X1 U2529 (.Y(n252), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1329]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN958_key_mem_1201_));
   AOI222X1 U2530 (.Y(n255), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[177]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[49]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1557_key_mem_305_));
   AOI222X1 U2531 (.Y(n254), 
	.C1(n2806), 
	.C0(key_mem[561]), 
	.B1(n2817), 
	.B0(key_mem[433]), 
	.A1(n2828), 
	.A0(FE_PHN1763_key_mem_689_));
   NAND4X1 U2532 (.Y(round_key[80]), 
	.D(n115), 
	.C(n114), 
	.B(n113), 
	.A(n112));
   AOI22X1 U2533 (.Y(n112), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1360]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN694_key_mem_1232_));
   AOI222X1 U2534 (.Y(n115), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[208]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[80]), 
	.A1(n21), 
	.A0(FE_PHN1493_key_mem_336_));
   AOI222X1 U2535 (.Y(n114), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[592]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[464]), 
	.A1(n2823), 
	.A0(FE_PHN1568_key_mem_720_));
   NAND4X1 U2536 (.Y(round_key[8]), 
	.D(n75), 
	.C(n74), 
	.B(n73), 
	.A(n72));
   AOI22X1 U2537 (.Y(n72), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1288]), 
	.A1(FE_OFN101_n30), 
	.A0(key_mem[1160]));
   AOI222X1 U2538 (.Y(n75), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[136]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[8]), 
	.A1(n21), 
	.A0(FE_PHN1632_key_mem_264_));
   AOI222X1 U2539 (.Y(n74), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[520]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[392]), 
	.A1(n2823), 
	.A0(FE_PHN1722_key_mem_648_));
   NAND4X1 U2540 (.Y(round_key[48]), 
	.D(n259), 
	.C(n258), 
	.B(n257), 
	.A(n256));
   AOI22X1 U2541 (.Y(n256), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1328]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN953_key_mem_1200_));
   AOI222X1 U2542 (.Y(n259), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[176]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[48]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1507_key_mem_304_));
   AOI222X1 U2543 (.Y(n258), 
	.C1(n2806), 
	.C0(key_mem[560]), 
	.B1(n2817), 
	.B0(key_mem[432]), 
	.A1(n2828), 
	.A0(FE_PHN1879_key_mem_688_));
   NAND4X1 U2544 (.Y(round_key[16]), 
	.D(n399), 
	.C(n398), 
	.B(n397), 
	.A(n396));
   AOI22X1 U2545 (.Y(n396), 
	.B1(n31), 
	.B0(key_mem[1296]), 
	.A1(n30), 
	.A0(key_mem[1168]));
   AOI222X1 U2546 (.Y(n399), 
	.C1(n23), 
	.C0(key_mem[144]), 
	.B1(n22), 
	.B0(key_mem[16]), 
	.A1(n21), 
	.A0(FE_PHN1672_key_mem_272_));
   AOI222X1 U2547 (.Y(n398), 
	.C1(n2806), 
	.C0(key_mem[528]), 
	.B1(n2818), 
	.B0(key_mem[400]), 
	.A1(n2823), 
	.A0(FE_PHN1657_key_mem_656_));
   NAND4X1 U2548 (.Y(round_key[112]), 
	.D(n483), 
	.C(n482), 
	.B(n481), 
	.A(n480));
   AOI22X1 U2549 (.Y(n480), 
	.B1(n31), 
	.B0(key_mem[1392]), 
	.A1(n30), 
	.A0(FE_PHN425_key_mem_1264_));
   AOI222X1 U2550 (.Y(n483), 
	.C1(n23), 
	.C0(key_mem[240]), 
	.B1(n22), 
	.B0(key_mem[112]), 
	.A1(n21), 
	.A0(FE_PHN1563_key_mem_368_));
   AOI222X1 U2551 (.Y(n482), 
	.C1(n2800), 
	.C0(key_mem[624]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[496]), 
	.A1(n2824), 
	.A0(FE_PHN1590_key_mem_752_));
   NAND4X1 U2552 (.Y(round_key[40]), 
	.D(n291), 
	.C(n290), 
	.B(n289), 
	.A(n288));
   AOI22X1 U2553 (.Y(n288), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1320]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN1005_key_mem_1192_));
   AOI222X1 U2554 (.Y(n291), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[168]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[40]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1562_key_mem_296_));
   AOI222X1 U2555 (.Y(n290), 
	.C1(n2806), 
	.C0(key_mem[552]), 
	.B1(n2817), 
	.B0(key_mem[424]), 
	.A1(n2828), 
	.A0(FE_PHN1696_key_mem_680_));
   NAND4X1 U2556 (.Y(round_key[104]), 
	.D(n519), 
	.C(n518), 
	.B(n517), 
	.A(n516));
   AOI22X1 U2557 (.Y(n516), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1384]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN432_key_mem_1256_));
   AOI222X1 U2558 (.Y(n519), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[232]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[104]), 
	.A1(n21), 
	.A0(FE_PHN1807_key_mem_360_));
   AOI222X1 U2559 (.Y(n518), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[616]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[488]), 
	.A1(n2823), 
	.A0(FE_PHN1550_key_mem_744_));
   NAND4X1 U2560 (.Y(round_key[23]), 
	.D(n367), 
	.C(n366), 
	.B(n365), 
	.A(n364));
   AOI22X1 U2561 (.Y(n364), 
	.B1(n31), 
	.B0(FE_PHN3094_key_mem_1303_), 
	.A1(n30), 
	.A0(FE_PHN585_key_mem_1175_));
   AOI222X1 U2562 (.Y(n367), 
	.C1(n23), 
	.C0(key_mem[151]), 
	.B1(n22), 
	.B0(key_mem[23]), 
	.A1(n21), 
	.A0(FE_PHN1715_key_mem_279_));
   AOI222X1 U2563 (.Y(n366), 
	.C1(n2800), 
	.C0(key_mem[535]), 
	.B1(FE_OFN99_n2811), 
	.B0(FE_PHN3209_key_mem_407_), 
	.A1(n2823), 
	.A0(FE_PHN1660_key_mem_663_));
   NAND4X1 U2564 (.Y(round_key[119]), 
	.D(n455), 
	.C(n454), 
	.B(n453), 
	.A(n452));
   AOI22X1 U2565 (.Y(n452), 
	.B1(n31), 
	.B0(key_mem[1399]), 
	.A1(n30), 
	.A0(FE_PHN984_key_mem_1271_));
   AOI222X1 U2566 (.Y(n455), 
	.C1(n23), 
	.C0(key_mem[247]), 
	.B1(n22), 
	.B0(key_mem[119]), 
	.A1(n21), 
	.A0(FE_PHN1598_key_mem_375_));
   AOI222X1 U2567 (.Y(n454), 
	.C1(n2800), 
	.C0(key_mem[631]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[503]), 
	.A1(n2824), 
	.A0(FE_PHN1723_key_mem_759_));
   NAND4X1 U2568 (.Y(round_key[87]), 
	.D(n87), 
	.C(n86), 
	.B(n85), 
	.A(n84));
   AOI22X1 U2569 (.Y(n84), 
	.B1(n31), 
	.B0(key_mem[1367]), 
	.A1(n30), 
	.A0(FE_PHN776_key_mem_1239_));
   AOI222X1 U2570 (.Y(n87), 
	.C1(n23), 
	.C0(key_mem[215]), 
	.B1(n22), 
	.B0(key_mem[87]), 
	.A1(n21), 
	.A0(FE_PHN1707_key_mem_343_));
   AOI222X1 U2571 (.Y(n86), 
	.C1(n2800), 
	.C0(key_mem[599]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[471]), 
	.A1(n2823), 
	.A0(key_mem[727]));
   NAND4X1 U2572 (.Y(round_key[55]), 
	.D(n227), 
	.C(n226), 
	.B(n225), 
	.A(n224));
   AOI22X1 U2573 (.Y(n224), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1335]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN1917_key_mem_1207_));
   AOI222X1 U2574 (.Y(n227), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[183]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[55]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1795_key_mem_311_));
   AOI222X1 U2575 (.Y(n226), 
	.C1(n2806), 
	.C0(key_mem[567]), 
	.B1(n2818), 
	.B0(key_mem[439]), 
	.A1(n2829), 
	.A0(FE_PHN939_key_mem_695_));
   NAND4X1 U2576 (.Y(round_key[71]), 
	.D(n155), 
	.C(n154), 
	.B(n153), 
	.A(n152));
   AOI22X1 U2577 (.Y(n152), 
	.B1(FE_OFN102_n31), 
	.B0(FE_PHN2828_key_mem_1351_), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN689_key_mem_1223_));
   AOI222X1 U2578 (.Y(n155), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[199]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[71]), 
	.A1(n21), 
	.A0(FE_PHN1543_key_mem_327_));
   AOI222X1 U2579 (.Y(n154), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[583]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[455]), 
	.A1(n2823), 
	.A0(FE_PHN1609_key_mem_711_));
   NAND4X1 U2580 (.Y(round_key[86]), 
	.D(n91), 
	.C(n90), 
	.B(n89), 
	.A(n88));
   AOI22X1 U2581 (.Y(n88), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1366]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN936_key_mem_1238_));
   AOI222X1 U2582 (.Y(n91), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[214]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[86]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1653_key_mem_342_));
   AOI222X1 U2583 (.Y(n90), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[598]), 
	.B1(n2817), 
	.B0(key_mem[470]), 
	.A1(n2823), 
	.A0(FE_PHN1646_key_mem_726_));
   NAND4X1 U2584 (.Y(round_key[54]), 
	.D(n231), 
	.C(n230), 
	.B(n229), 
	.A(n228));
   AOI22X1 U2585 (.Y(n228), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1334]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN1021_key_mem_1206_));
   AOI222X1 U2586 (.Y(n231), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[182]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[54]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1547_key_mem_310_));
   AOI222X1 U2587 (.Y(n230), 
	.C1(n2806), 
	.C0(key_mem[566]), 
	.B1(n2818), 
	.B0(key_mem[438]), 
	.A1(n2829), 
	.A0(FE_PHN1779_key_mem_694_));
   NAND4X1 U2588 (.Y(round_key[22]), 
	.D(n371), 
	.C(n370), 
	.B(n369), 
	.A(n368));
   AOI22X1 U2589 (.Y(n368), 
	.B1(n31), 
	.B0(FE_PHN2835_key_mem_1302_), 
	.A1(n30), 
	.A0(FE_PHN1000_key_mem_1174_));
   AOI222X1 U2590 (.Y(n371), 
	.C1(n23), 
	.C0(key_mem[150]), 
	.B1(n22), 
	.B0(key_mem[22]), 
	.A1(n21), 
	.A0(FE_PHN1622_key_mem_278_));
   AOI222X1 U2591 (.Y(n370), 
	.C1(n2800), 
	.C0(key_mem[534]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[406]), 
	.A1(n2823), 
	.A0(FE_PHN1687_key_mem_662_));
   NAND4X1 U2592 (.Y(round_key[118]), 
	.D(n459), 
	.C(n458), 
	.B(n457), 
	.A(n456));
   AOI22X1 U2593 (.Y(n456), 
	.B1(n31), 
	.B0(key_mem[1398]), 
	.A1(n30), 
	.A0(FE_PHN990_key_mem_1270_));
   AOI222X1 U2594 (.Y(n459), 
	.C1(n23), 
	.C0(key_mem[246]), 
	.B1(n22), 
	.B0(key_mem[118]), 
	.A1(n21), 
	.A0(FE_PHN1726_key_mem_374_));
   AOI222X1 U2595 (.Y(n458), 
	.C1(n2800), 
	.C0(key_mem[630]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[502]), 
	.A1(n2824), 
	.A0(FE_PHN1751_key_mem_758_));
   NAND4X1 U2596 (.Y(round_key[85]), 
	.D(n95), 
	.C(n94), 
	.B(n93), 
	.A(n92));
   AOI22X1 U2597 (.Y(n92), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1365]), 
	.A1(FE_OFN101_n30), 
	.A0(key_mem[1237]));
   AOI222X1 U2598 (.Y(n95), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[213]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[85]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1714_key_mem_341_));
   AOI222X1 U2599 (.Y(n94), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[597]), 
	.B1(n2817), 
	.B0(key_mem[469]), 
	.A1(n2823), 
	.A0(FE_PHN1556_key_mem_725_));
   NAND4X1 U2600 (.Y(round_key[53]), 
	.D(n235), 
	.C(n234), 
	.B(n233), 
	.A(n232));
   AOI22X1 U2601 (.Y(n232), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1333]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN1024_key_mem_1205_));
   AOI222X1 U2602 (.Y(n235), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[181]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[53]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1717_key_mem_309_));
   AOI222X1 U2603 (.Y(n234), 
	.C1(n2806), 
	.C0(key_mem[565]), 
	.B1(n2818), 
	.B0(key_mem[437]), 
	.A1(n2829), 
	.A0(FE_PHN1731_key_mem_693_));
   NAND4X1 U2604 (.Y(round_key[21]), 
	.D(n375), 
	.C(n374), 
	.B(n373), 
	.A(n372));
   AOI22X1 U2605 (.Y(n372), 
	.B1(n31), 
	.B0(key_mem[1301]), 
	.A1(n30), 
	.A0(FE_PHN768_key_mem_1173_));
   AOI222X1 U2606 (.Y(n375), 
	.C1(n23), 
	.C0(key_mem[149]), 
	.B1(n22), 
	.B0(key_mem[21]), 
	.A1(n21), 
	.A0(FE_PHN1484_key_mem_277_));
   AOI222X1 U2607 (.Y(n374), 
	.C1(n2800), 
	.C0(key_mem[533]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[405]), 
	.A1(n2823), 
	.A0(FE_PHN1797_key_mem_661_));
   NAND4X1 U2608 (.Y(round_key[77]), 
	.D(n131), 
	.C(n130), 
	.B(n129), 
	.A(n128));
   AOI22X1 U2609 (.Y(n128), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1357]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN934_key_mem_1229_));
   AOI222X1 U2610 (.Y(n131), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[205]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[77]), 
	.A1(n21), 
	.A0(FE_PHN1472_key_mem_333_));
   AOI222X1 U2611 (.Y(n130), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[589]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[461]), 
	.A1(n2823), 
	.A0(FE_PHN1523_key_mem_717_));
   NAND4X1 U2612 (.Y(round_key[52]), 
	.D(n239), 
	.C(n238), 
	.B(n237), 
	.A(n236));
   AOI22X1 U2613 (.Y(n236), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1332]), 
	.A1(FE_OFN101_n30), 
	.A0(key_mem[1204]));
   AOI222X1 U2614 (.Y(n239), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[180]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[52]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1691_key_mem_308_));
   AOI222X1 U2615 (.Y(n238), 
	.C1(n2806), 
	.C0(key_mem[564]), 
	.B1(n2818), 
	.B0(key_mem[436]), 
	.A1(n2829), 
	.A0(FE_PHN1638_key_mem_692_));
   NAND4X1 U2616 (.Y(round_key[19]), 
	.D(n387), 
	.C(n386), 
	.B(n385), 
	.A(n384));
   AOI22X1 U2617 (.Y(n384), 
	.B1(n31), 
	.B0(FE_PHN3435_key_mem_1299_), 
	.A1(n30), 
	.A0(FE_PHN2839_key_mem_1171_));
   AOI222X1 U2618 (.Y(n387), 
	.C1(n23), 
	.C0(key_mem[147]), 
	.B1(n22), 
	.B0(FE_PHN3188_key_mem_19_), 
	.A1(n21), 
	.A0(FE_PHN763_key_mem_275_));
   AOI222X1 U2619 (.Y(n386), 
	.C1(n2800), 
	.C0(key_mem[531]), 
	.B1(FE_OFN99_n2811), 
	.B0(FE_PHN3218_key_mem_403_), 
	.A1(n2823), 
	.A0(FE_PHN1744_key_mem_659_));
   NAND4X1 U2620 (.Y(round_key[75]), 
	.D(n139), 
	.C(n138), 
	.B(n137), 
	.A(n136));
   AOI22X1 U2621 (.Y(n136), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1355]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN975_key_mem_1227_));
   AOI222X1 U2622 (.Y(n139), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[203]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[75]), 
	.A1(n21), 
	.A0(FE_PHN1475_key_mem_331_));
   AOI222X1 U2623 (.Y(n138), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[587]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[459]), 
	.A1(n2823), 
	.A0(FE_PHN1678_key_mem_715_));
   NAND4X1 U2624 (.Y(round_key[1]), 
	.D(n383), 
	.C(n382), 
	.B(n381), 
	.A(n380));
   AOI22X1 U2625 (.Y(n380), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1281]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN1883_key_mem_1153_));
   AOI222X1 U2626 (.Y(n383), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[129]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[1]), 
	.A1(n21), 
	.A0(FE_PHN1553_key_mem_257_));
   AOI222X1 U2627 (.Y(n382), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[513]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[385]), 
	.A1(n2823), 
	.A0(FE_PHN683_key_mem_641_));
   NAND4X1 U2628 (.Y(round_key[32]), 
	.D(n327), 
	.C(n326), 
	.B(n325), 
	.A(n324));
   AOI22X1 U2629 (.Y(n324), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1312]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN426_key_mem_1184_));
   AOI222X1 U2630 (.Y(n327), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[160]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[32]), 
	.A1(n21), 
	.A0(FE_PHN1684_key_mem_288_));
   AOI222X1 U2631 (.Y(n326), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[544]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[416]), 
	.A1(n2827), 
	.A0(FE_PHN1581_key_mem_672_));
   NAND4X1 U2632 (.Y(round_key[20]), 
	.D(n379), 
	.C(n378), 
	.B(n377), 
	.A(n376));
   AOI22X1 U2633 (.Y(n376), 
	.B1(n31), 
	.B0(key_mem[1300]), 
	.A1(n30), 
	.A0(FE_PHN698_key_mem_1172_));
   AOI222X1 U2634 (.Y(n379), 
	.C1(n23), 
	.C0(key_mem[148]), 
	.B1(n22), 
	.B0(key_mem[20]), 
	.A1(n21), 
	.A0(FE_PHN1522_key_mem_276_));
   AOI222X1 U2635 (.Y(n378), 
	.C1(n2800), 
	.C0(key_mem[532]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[404]), 
	.A1(n2823), 
	.A0(FE_PHN1724_key_mem_660_));
   NAND4X1 U2636 (.Y(round_key[116]), 
	.D(n467), 
	.C(n466), 
	.B(n465), 
	.A(n464));
   AOI22X1 U2637 (.Y(n464), 
	.B1(n31), 
	.B0(key_mem[1396]), 
	.A1(n30), 
	.A0(FE_PHN935_key_mem_1268_));
   AOI222X1 U2638 (.Y(n467), 
	.C1(n23), 
	.C0(key_mem[244]), 
	.B1(n22), 
	.B0(key_mem[116]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1580_key_mem_372_));
   AOI222X1 U2639 (.Y(n466), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[628]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[500]), 
	.A1(n2824), 
	.A0(FE_PHN1631_key_mem_756_));
   NAND4X1 U2640 (.Y(round_key[83]), 
	.D(n103), 
	.C(n102), 
	.B(n101), 
	.A(n100));
   AOI22X1 U2641 (.Y(n100), 
	.B1(n31), 
	.B0(key_mem[1363]), 
	.A1(n30), 
	.A0(FE_PHN972_key_mem_1235_));
   AOI222X1 U2642 (.Y(n103), 
	.C1(n23), 
	.C0(key_mem[211]), 
	.B1(n22), 
	.B0(key_mem[83]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1464_key_mem_339_));
   AOI222X1 U2643 (.Y(n102), 
	.C1(n2800), 
	.C0(key_mem[595]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[467]), 
	.A1(n2823), 
	.A0(FE_PHN1770_key_mem_723_));
   NAND4X1 U2644 (.Y(round_key[7]), 
	.D(n119), 
	.C(n118), 
	.B(n117), 
	.A(n116));
   AOI22X1 U2645 (.Y(n116), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1287]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN584_key_mem_1159_));
   AOI222X1 U2646 (.Y(n119), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[135]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[7]), 
	.A1(n21), 
	.A0(FE_PHN1682_key_mem_263_));
   AOI222X1 U2647 (.Y(n118), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[519]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[391]), 
	.A1(n2823), 
	.A0(FE_PHN1848_key_mem_647_));
   NAND4X1 U2648 (.Y(round_key[79]), 
	.D(n123), 
	.C(n122), 
	.B(n121), 
	.A(n120));
   AOI22X1 U2649 (.Y(n120), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1359]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN949_key_mem_1231_));
   AOI222X1 U2650 (.Y(n123), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[207]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[79]), 
	.A1(n21), 
	.A0(FE_PHN1494_key_mem_335_));
   AOI222X1 U2651 (.Y(n122), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[591]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[463]), 
	.A1(n2823), 
	.A0(FE_PHN1530_key_mem_719_));
   NAND4X1 U2652 (.Y(round_key[14]), 
	.D(n407), 
	.C(n406), 
	.B(n405), 
	.A(n404));
   AOI22X1 U2653 (.Y(n404), 
	.B1(n31), 
	.B0(key_mem[1294]), 
	.A1(n30), 
	.A0(FE_PHN798_key_mem_1166_));
   AOI222X1 U2654 (.Y(n407), 
	.C1(n23), 
	.C0(key_mem[142]), 
	.B1(n22), 
	.B0(key_mem[14]), 
	.A1(n21), 
	.A0(FE_PHN1626_key_mem_270_));
   AOI222X1 U2655 (.Y(n406), 
	.C1(n2806), 
	.C0(key_mem[526]), 
	.B1(n2818), 
	.B0(key_mem[398]), 
	.A1(n2823), 
	.A0(FE_PHN1577_key_mem_654_));
   NAND4X1 U2656 (.Y(round_key[117]), 
	.D(n463), 
	.C(n462), 
	.B(n461), 
	.A(n460));
   AOI22X1 U2657 (.Y(n460), 
	.B1(n31), 
	.B0(key_mem[1397]), 
	.A1(n30), 
	.A0(key_mem[1269]));
   AOI222X1 U2658 (.Y(n463), 
	.C1(n23), 
	.C0(key_mem[245]), 
	.B1(n22), 
	.B0(key_mem[117]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1498_key_mem_373_));
   AOI222X1 U2659 (.Y(n462), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[629]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[501]), 
	.A1(n2824), 
	.A0(FE_PHN1679_key_mem_757_));
   NAND4X1 U2660 (.Y(round_key[44]), 
	.D(n275), 
	.C(n274), 
	.B(n273), 
	.A(n272));
   AOI22X1 U2661 (.Y(n272), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1324]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN929_key_mem_1196_));
   AOI222X1 U2662 (.Y(n275), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[172]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[44]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1544_key_mem_300_));
   AOI222X1 U2663 (.Y(n274), 
	.C1(n2806), 
	.C0(key_mem[556]), 
	.B1(n2817), 
	.B0(key_mem[428]), 
	.A1(n2828), 
	.A0(FE_PHN1776_key_mem_684_));
   NAND4X1 U2664 (.Y(round_key[67]), 
	.D(n175), 
	.C(n174), 
	.B(n173), 
	.A(n172));
   AOI22X1 U2665 (.Y(n172), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1347]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN1006_key_mem_1219_));
   AOI222X1 U2666 (.Y(n175), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[195]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[67]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1683_key_mem_323_));
   AOI222X1 U2667 (.Y(n174), 
	.C1(n2800), 
	.C0(key_mem[579]), 
	.B1(n2818), 
	.B0(key_mem[451]), 
	.A1(n2828), 
	.A0(FE_PHN1750_key_mem_707_));
   NAND4X1 U2668 (.Y(round_key[11]), 
	.D(n451), 
	.C(n450), 
	.B(n449), 
	.A(n448));
   AOI22X1 U2669 (.Y(n448), 
	.B1(n31), 
	.B0(key_mem[1291]), 
	.A1(n30), 
	.A0(FE_PHN974_key_mem_1163_));
   AOI222X1 U2670 (.Y(n451), 
	.C1(n23), 
	.C0(key_mem[139]), 
	.B1(n22), 
	.B0(key_mem[11]), 
	.A1(n21), 
	.A0(key_mem[267]));
   AOI222X1 U2671 (.Y(n450), 
	.C1(n2800), 
	.C0(key_mem[523]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[395]), 
	.A1(n2824), 
	.A0(key_mem[651]));
   NAND4X1 U2672 (.Y(round_key[74]), 
	.D(n143), 
	.C(n142), 
	.B(n141), 
	.A(n140));
   AOI22X1 U2673 (.Y(n140), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1354]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN692_key_mem_1226_));
   AOI222X1 U2674 (.Y(n143), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[202]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[74]), 
	.A1(n21), 
	.A0(FE_PHN1603_key_mem_330_));
   AOI222X1 U2675 (.Y(n142), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[586]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[458]), 
	.A1(n2823), 
	.A0(FE_PHN1495_key_mem_714_));
   NAND4X1 U2676 (.Y(round_key[72]), 
	.D(n151), 
	.C(n150), 
	.B(n149), 
	.A(n148));
   AOI22X1 U2677 (.Y(n148), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1352]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN431_key_mem_1224_));
   AOI222X1 U2678 (.Y(n151), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[200]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[72]), 
	.A1(n21), 
	.A0(FE_PHN1742_key_mem_328_));
   AOI222X1 U2679 (.Y(n150), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[584]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[456]), 
	.A1(n2823), 
	.A0(FE_PHN1524_key_mem_712_));
   NAND4X1 U2680 (.Y(round_key[15]), 
	.D(n403), 
	.C(n402), 
	.B(n401), 
	.A(n400));
   AOI22X1 U2681 (.Y(n400), 
	.B1(n31), 
	.B0(FE_PHN2840_key_mem_1295_), 
	.A1(n30), 
	.A0(FE_PHN430_key_mem_1167_));
   AOI222X1 U2682 (.Y(n403), 
	.C1(n23), 
	.C0(FE_PHN3420_key_mem_143_), 
	.B1(n22), 
	.B0(FE_PHN3283_key_mem_15_), 
	.A1(n21), 
	.A0(FE_PHN1504_key_mem_271_));
   AOI222X1 U2683 (.Y(n402), 
	.C1(n2806), 
	.C0(key_mem[527]), 
	.B1(n2818), 
	.B0(FE_PHN3204_key_mem_399_), 
	.A1(n2823), 
	.A0(FE_PHN1588_key_mem_655_));
   NAND4X1 U2684 (.Y(round_key[78]), 
	.D(n127), 
	.C(n126), 
	.B(n125), 
	.A(n124));
   AOI22X1 U2685 (.Y(n124), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1358]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN591_key_mem_1230_));
   AOI222X1 U2686 (.Y(n127), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[206]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[78]), 
	.A1(n21), 
	.A0(FE_PHN1826_key_mem_334_));
   AOI222X1 U2687 (.Y(n126), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[590]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[462]), 
	.A1(n2823), 
	.A0(FE_PHN1521_key_mem_718_));
   NAND4X1 U2688 (.Y(round_key[13]), 
	.D(n411), 
	.C(n410), 
	.B(n409), 
	.A(n408));
   AOI22X1 U2689 (.Y(n408), 
	.B1(n31), 
	.B0(key_mem[1293]), 
	.A1(n30), 
	.A0(key_mem[1165]));
   AOI222X1 U2690 (.Y(n411), 
	.C1(n23), 
	.C0(key_mem[141]), 
	.B1(n22), 
	.B0(key_mem[13]), 
	.A1(n21), 
	.A0(FE_PHN1727_key_mem_269_));
   AOI222X1 U2691 (.Y(n410), 
	.C1(n2806), 
	.C0(key_mem[525]), 
	.B1(n2818), 
	.B0(key_mem[397]), 
	.A1(n2823), 
	.A0(key_mem[653]));
   NAND4X1 U2692 (.Y(round_key[76]), 
	.D(n135), 
	.C(n134), 
	.B(n133), 
	.A(n132));
   AOI22X1 U2693 (.Y(n132), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1356]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN960_key_mem_1228_));
   AOI222X1 U2694 (.Y(n135), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[204]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[76]), 
	.A1(n21), 
	.A0(FE_PHN1514_key_mem_332_));
   AOI222X1 U2695 (.Y(n134), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[588]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[460]), 
	.A1(n2823), 
	.A0(FE_PHN1695_key_mem_716_));
   NAND4X1 U2696 (.Y(round_key[100]), 
	.D(n535), 
	.C(n534), 
	.B(n533), 
	.A(n532));
   AOI22X1 U2697 (.Y(n532), 
	.B1(n31), 
	.B0(key_mem[1380]), 
	.A1(n30), 
	.A0(FE_PHN688_key_mem_1252_));
   AOI222X1 U2698 (.Y(n535), 
	.C1(n23), 
	.C0(key_mem[228]), 
	.B1(n22), 
	.B0(key_mem[100]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1549_key_mem_356_));
   AOI222X1 U2699 (.Y(n534), 
	.C1(n2800), 
	.C0(key_mem[612]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[484]), 
	.A1(n2823), 
	.A0(key_mem[740]));
   NAND4X1 U2700 (.Y(round_key[84]), 
	.D(n99), 
	.C(n98), 
	.B(n97), 
	.A(n96));
   AOI22X1 U2701 (.Y(n96), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1364]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN968_key_mem_1236_));
   AOI222X1 U2702 (.Y(n99), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[212]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[84]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1620_key_mem_340_));
   AOI222X1 U2703 (.Y(n98), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[596]), 
	.B1(n2817), 
	.B0(key_mem[468]), 
	.A1(n2823), 
	.A0(FE_PHN1831_key_mem_724_));
   NAND4X1 U2704 (.Y(round_key[51]), 
	.D(n243), 
	.C(n242), 
	.B(n241), 
	.A(n240));
   AOI22X1 U2705 (.Y(n240), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1331]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN942_key_mem_1203_));
   AOI222X1 U2706 (.Y(n243), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[179]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[51]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1633_key_mem_307_));
   AOI222X1 U2707 (.Y(n242), 
	.C1(n2806), 
	.C0(key_mem[563]), 
	.B1(n2818), 
	.B0(key_mem[435]), 
	.A1(n2829), 
	.A0(FE_PHN1476_key_mem_691_));
   NAND4X1 U2708 (.Y(round_key[106]), 
	.D(n511), 
	.C(n510), 
	.B(n509), 
	.A(n508));
   AOI22X1 U2709 (.Y(n508), 
	.B1(n31), 
	.B0(FE_PHN2810_key_mem_1386_), 
	.A1(n30), 
	.A0(FE_PHN427_key_mem_1258_));
   AOI222X1 U2710 (.Y(n511), 
	.C1(n23), 
	.C0(FE_PHN3423_key_mem_234_), 
	.B1(n22), 
	.B0(FE_PHN3185_key_mem_106_), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1594_key_mem_362_));
   AOI222X1 U2711 (.Y(n510), 
	.C1(n2800), 
	.C0(FE_PHN3415_key_mem_618_), 
	.B1(FE_OFN99_n2811), 
	.B0(FE_PHN3422_key_mem_490_), 
	.A1(n2823), 
	.A0(FE_PHN3215_key_mem_746_));
   NAND4X1 U2712 (.Y(round_key[41]), 
	.D(n287), 
	.C(n286), 
	.B(n285), 
	.A(n284));
   AOI22X1 U2713 (.Y(n284), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1321]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN1029_key_mem_1193_));
   AOI222X1 U2714 (.Y(n287), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[169]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[41]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1729_key_mem_297_));
   AOI222X1 U2715 (.Y(n286), 
	.C1(n2806), 
	.C0(key_mem[553]), 
	.B1(n2817), 
	.B0(key_mem[425]), 
	.A1(n2828), 
	.A0(FE_PHN1564_key_mem_681_));
   NAND4X1 U2716 (.Y(round_key[64]), 
	.D(n187), 
	.C(n186), 
	.B(n185), 
	.A(n184));
   AOI22X1 U2717 (.Y(n184), 
	.B1(FE_OFN102_n31), 
	.B0(FE_PHN969_key_mem_1344_), 
	.A1(FE_OFN101_n30), 
	.A0(key_mem[1216]));
   AOI222X1 U2718 (.Y(n187), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[192]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[64]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1555_key_mem_320_));
   AOI222X1 U2719 (.Y(n186), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[576]), 
	.B1(n2818), 
	.B0(key_mem[448]), 
	.A1(n2828), 
	.A0(FE_PHN1721_key_mem_704_));
   NAND4X1 U2720 (.Y(round_key[103]), 
	.D(n523), 
	.C(n522), 
	.B(n521), 
	.A(n520));
   AOI22X1 U2721 (.Y(n520), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1383]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN1877_key_mem_1255_));
   AOI222X1 U2722 (.Y(n523), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[231]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[103]), 
	.A1(n21), 
	.A0(FE_PHN1757_key_mem_359_));
   AOI222X1 U2723 (.Y(n522), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[615]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[487]), 
	.A1(n2823), 
	.A0(FE_PHN580_key_mem_743_));
   NAND4X1 U2724 (.Y(round_key[47]), 
	.D(n263), 
	.C(n262), 
	.B(n261), 
	.A(n260));
   AOI22X1 U2725 (.Y(n260), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1327]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN1008_key_mem_1199_));
   AOI222X1 U2726 (.Y(n263), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[175]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[47]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1600_key_mem_303_));
   AOI222X1 U2727 (.Y(n262), 
	.C1(n2806), 
	.C0(key_mem[559]), 
	.B1(n2817), 
	.B0(key_mem[431]), 
	.A1(n2828), 
	.A0(FE_PHN1663_key_mem_687_));
   NAND4X1 U2728 (.Y(round_key[70]), 
	.D(n159), 
	.C(n158), 
	.B(n157), 
	.A(n156));
   AOI22X1 U2729 (.Y(n156), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1350]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN1010_key_mem_1222_));
   AOI222X1 U2730 (.Y(n159), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[198]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[70]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1479_key_mem_326_));
   AOI222X1 U2731 (.Y(n158), 
	.C1(n2800), 
	.C0(key_mem[582]), 
	.B1(n2818), 
	.B0(key_mem[454]), 
	.A1(n2828), 
	.A0(FE_PHN1702_key_mem_710_));
   NAND4X1 U2732 (.Y(round_key[102]), 
	.D(n527), 
	.C(n526), 
	.B(n525), 
	.A(n524));
   AOI22X1 U2733 (.Y(n524), 
	.B1(FE_OFN102_n31), 
	.B0(FE_PHN2836_key_mem_1382_), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN699_key_mem_1254_));
   AOI222X1 U2734 (.Y(n527), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[230]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[102]), 
	.A1(n21), 
	.A0(FE_PHN1655_key_mem_358_));
   AOI222X1 U2735 (.Y(n526), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[614]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[486]), 
	.A1(n2823), 
	.A0(FE_PHN1668_key_mem_742_));
   NAND4X1 U2736 (.Y(round_key[46]), 
	.D(n267), 
	.C(n266), 
	.B(n265), 
	.A(n264));
   AOI22X1 U2737 (.Y(n264), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1326]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN955_key_mem_1198_));
   AOI222X1 U2738 (.Y(n267), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[174]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[46]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1785_key_mem_302_));
   AOI222X1 U2739 (.Y(n266), 
	.C1(n2806), 
	.C0(key_mem[558]), 
	.B1(n2817), 
	.B0(key_mem[430]), 
	.A1(n2828), 
	.A0(FE_PHN1593_key_mem_686_));
   NAND4X1 U2740 (.Y(round_key[69]), 
	.D(n167), 
	.C(n166), 
	.B(n165), 
	.A(n164));
   AOI22X1 U2741 (.Y(n164), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1349]), 
	.A1(FE_OFN101_n30), 
	.A0(key_mem[1221]));
   AOI222X1 U2742 (.Y(n167), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[197]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[69]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1689_key_mem_325_));
   AOI222X1 U2743 (.Y(n166), 
	.C1(n2800), 
	.C0(key_mem[581]), 
	.B1(n2818), 
	.B0(key_mem[453]), 
	.A1(n2828), 
	.A0(FE_PHN1794_key_mem_709_));
   NAND4X1 U2744 (.Y(round_key[101]), 
	.D(n531), 
	.C(n530), 
	.B(n529), 
	.A(n528));
   AOI22X1 U2745 (.Y(n528), 
	.B1(n31), 
	.B0(key_mem[1381]), 
	.A1(n30), 
	.A0(FE_PHN1014_key_mem_1253_));
   AOI222X1 U2746 (.Y(n531), 
	.C1(n23), 
	.C0(key_mem[229]), 
	.B1(n22), 
	.B0(key_mem[101]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1583_key_mem_357_));
   AOI222X1 U2747 (.Y(n530), 
	.C1(n2800), 
	.C0(key_mem[613]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[485]), 
	.A1(n2823), 
	.A0(FE_PHN1606_key_mem_741_));
   NAND4X1 U2748 (.Y(round_key[45]), 
	.D(n271), 
	.C(n270), 
	.B(n269), 
	.A(n268));
   AOI22X1 U2749 (.Y(n268), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1325]), 
	.A1(FE_OFN101_n30), 
	.A0(key_mem[1197]));
   AOI222X1 U2750 (.Y(n271), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[173]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[45]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1650_key_mem_301_));
   AOI222X1 U2751 (.Y(n270), 
	.C1(n2806), 
	.C0(key_mem[557]), 
	.B1(n2817), 
	.B0(key_mem[429]), 
	.A1(n2828), 
	.A0(FE_PHN1630_key_mem_685_));
   NAND4X1 U2752 (.Y(round_key[68]), 
	.D(n171), 
	.C(n170), 
	.B(n169), 
	.A(n168));
   AOI22X1 U2753 (.Y(n168), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1348]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN977_key_mem_1220_));
   AOI222X1 U2754 (.Y(n171), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[196]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[68]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1716_key_mem_324_));
   AOI222X1 U2755 (.Y(n170), 
	.C1(n2800), 
	.C0(key_mem[580]), 
	.B1(n2818), 
	.B0(key_mem[452]), 
	.A1(n2828), 
	.A0(FE_PHN1755_key_mem_708_));
   NAND4X1 U2756 (.Y(round_key[12]), 
	.D(n415), 
	.C(n414), 
	.B(n413), 
	.A(n412));
   AOI22X1 U2757 (.Y(n412), 
	.B1(n31), 
	.B0(key_mem[1292]), 
	.A1(n30), 
	.A0(key_mem[1164]));
   AOI222X1 U2758 (.Y(n415), 
	.C1(n23), 
	.C0(key_mem[140]), 
	.B1(n22), 
	.B0(key_mem[12]), 
	.A1(n21), 
	.A0(FE_PHN1571_key_mem_268_));
   AOI222X1 U2759 (.Y(n414), 
	.C1(n2806), 
	.C0(key_mem[524]), 
	.B1(n2818), 
	.B0(key_mem[396]), 
	.A1(n2823), 
	.A0(FE_PHN914_key_mem_652_));
   NAND4X1 U2760 (.Y(round_key[36]), 
	.D(n311), 
	.C(n310), 
	.B(n309), 
	.A(n308));
   AOI22X1 U2761 (.Y(n308), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1316]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN1720_key_mem_1188_));
   AOI222X1 U2762 (.Y(n311), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[164]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[36]), 
	.A1(n21), 
	.A0(FE_PHN1525_key_mem_292_));
   AOI222X1 U2763 (.Y(n310), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[548]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[420]), 
	.A1(n2827), 
	.A0(FE_PHN917_key_mem_676_));
   NAND4X1 U2764 (.Y(round_key[108]), 
	.D(n503), 
	.C(n502), 
	.B(n501), 
	.A(n500));
   AOI22X1 U2765 (.Y(n500), 
	.B1(n31), 
	.B0(key_mem[1388]), 
	.A1(n30), 
	.A0(FE_PHN947_key_mem_1260_));
   AOI222X1 U2766 (.Y(n503), 
	.C1(n23), 
	.C0(key_mem[236]), 
	.B1(n22), 
	.B0(key_mem[108]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1607_key_mem_364_));
   AOI222X1 U2767 (.Y(n502), 
	.C1(n2800), 
	.C0(key_mem[620]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[492]), 
	.A1(n2823), 
	.A0(FE_PHN1473_key_mem_748_));
   NAND4X1 U2768 (.Y(round_key[43]), 
	.D(n279), 
	.C(n278), 
	.B(n277), 
	.A(n276));
   AOI22X1 U2769 (.Y(n276), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1323]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN943_key_mem_1195_));
   AOI222X1 U2770 (.Y(n279), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[171]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[43]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1545_key_mem_299_));
   AOI222X1 U2771 (.Y(n278), 
	.C1(n2806), 
	.C0(key_mem[555]), 
	.B1(n2817), 
	.B0(key_mem[427]), 
	.A1(n2828), 
	.A0(FE_PHN1575_key_mem_683_));
   NAND4X1 U2772 (.Y(round_key[66]), 
	.D(n179), 
	.C(n178), 
	.B(n177), 
	.A(n176));
   AOI22X1 U2773 (.Y(n176), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1346]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN785_key_mem_1218_));
   AOI222X1 U2774 (.Y(n179), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[194]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[66]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1667_key_mem_322_));
   AOI222X1 U2775 (.Y(n178), 
	.C1(n2800), 
	.C0(key_mem[578]), 
	.B1(n2818), 
	.B0(key_mem[450]), 
	.A1(n2828), 
	.A0(FE_PHN1561_key_mem_706_));
   NAND4X1 U2776 (.Y(round_key[0]), 
	.D(n539), 
	.C(n538), 
	.B(n537), 
	.A(n536));
   AOI22X1 U2777 (.Y(n536), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1280]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN1734_key_mem_1152_));
   AOI222X1 U2778 (.Y(n539), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[128]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[0]), 
	.A1(n21), 
	.A0(FE_PHN1711_key_mem_256_));
   AOI222X1 U2779 (.Y(n538), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[512]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[384]), 
	.A1(n2823), 
	.A0(FE_PHN684_key_mem_640_));
   NAND4X1 U2780 (.Y(round_key[39]), 
	.D(n299), 
	.C(n298), 
	.B(n297), 
	.A(n296));
   AOI22X1 U2781 (.Y(n296), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1319]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN1800_key_mem_1191_));
   AOI222X1 U2782 (.Y(n299), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[167]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[39]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1511_key_mem_295_));
   AOI222X1 U2783 (.Y(n298), 
	.C1(n2806), 
	.C0(key_mem[551]), 
	.B1(n2817), 
	.B0(key_mem[423]), 
	.A1(n2828), 
	.A0(FE_PHN1565_key_mem_679_));
   NAND4X1 U2784 (.Y(round_key[111]), 
	.D(n487), 
	.C(n486), 
	.B(n485), 
	.A(n484));
   AOI22X1 U2785 (.Y(n484), 
	.B1(n31), 
	.B0(FE_PHN3419_key_mem_1391_), 
	.A1(n30), 
	.A0(FE_PHN2842_key_mem_1263_));
   AOI222X1 U2786 (.Y(n487), 
	.C1(n23), 
	.C0(FE_PHN3427_key_mem_239_), 
	.B1(n22), 
	.B0(FE_PHN3187_key_mem_111_), 
	.A1(n21), 
	.A0(FE_PHN424_key_mem_367_));
   AOI222X1 U2787 (.Y(n486), 
	.C1(n2800), 
	.C0(FE_PHN3413_key_mem_623_), 
	.B1(FE_OFN99_n2811), 
	.B0(FE_PHN3213_key_mem_495_), 
	.A1(n2824), 
	.A0(FE_PHN1613_key_mem_751_));
   NAND4X1 U2788 (.Y(round_key[6]), 
	.D(n163), 
	.C(n162), 
	.B(n161), 
	.A(n160));
   AOI22X1 U2789 (.Y(n160), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1286]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN980_key_mem_1158_));
   AOI222X1 U2790 (.Y(n163), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[134]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[6]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1699_key_mem_262_));
   AOI222X1 U2791 (.Y(n162), 
	.C1(n2800), 
	.C0(key_mem[518]), 
	.B1(n2818), 
	.B0(key_mem[390]), 
	.A1(n2828), 
	.A0(key_mem[646]));
   NAND4X1 U2792 (.Y(round_key[38]), 
	.D(n303), 
	.C(n302), 
	.B(n301), 
	.A(n300));
   AOI22X1 U2793 (.Y(n300), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1318]), 
	.A1(FE_OFN101_n30), 
	.A0(key_mem[1190]));
   AOI222X1 U2794 (.Y(n303), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[166]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[38]), 
	.A1(n21), 
	.A0(FE_PHN1601_key_mem_294_));
   AOI222X1 U2795 (.Y(n302), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[550]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[422]), 
	.A1(n2827), 
	.A0(FE_PHN1579_key_mem_678_));
   NAND4X1 U2796 (.Y(round_key[110]), 
	.D(n491), 
	.C(n490), 
	.B(n489), 
	.A(n488));
   AOI22X1 U2797 (.Y(n488), 
	.B1(n31), 
	.B0(FE_PHN592_key_mem_1390_), 
	.A1(n30), 
	.A0(FE_PHN2831_key_mem_1262_));
   AOI222X1 U2798 (.Y(n491), 
	.C1(n23), 
	.C0(key_mem[238]), 
	.B1(n22), 
	.B0(key_mem[110]), 
	.A1(n21), 
	.A0(FE_PHN1538_key_mem_366_));
   AOI222X1 U2799 (.Y(n490), 
	.C1(n2800), 
	.C0(key_mem[622]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[494]), 
	.A1(n2824), 
	.A0(FE_PHN1636_key_mem_750_));
   NAND4X1 U2800 (.Y(round_key[5]), 
	.D(n207), 
	.C(n206), 
	.B(n205), 
	.A(n204));
   AOI22X1 U2801 (.Y(n204), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1285]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN989_key_mem_1157_));
   AOI222X1 U2802 (.Y(n207), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[133]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[5]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1652_key_mem_261_));
   AOI222X1 U2803 (.Y(n206), 
	.C1(n2806), 
	.C0(key_mem[517]), 
	.B1(n2818), 
	.B0(key_mem[389]), 
	.A1(n2829), 
	.A0(FE_PHN1624_key_mem_645_));
   NAND4X1 U2804 (.Y(round_key[37]), 
	.D(n307), 
	.C(n306), 
	.B(n305), 
	.A(n304));
   AOI22X1 U2805 (.Y(n304), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1317]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN1083_key_mem_1189_));
   AOI222X1 U2806 (.Y(n307), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[165]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[37]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1616_key_mem_293_));
   AOI222X1 U2807 (.Y(n306), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[549]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[421]), 
	.A1(n2827), 
	.A0(FE_PHN1661_key_mem_677_));
   NAND4X1 U2808 (.Y(round_key[109]), 
	.D(n499), 
	.C(n498), 
	.B(n497), 
	.A(n496));
   AOI22X1 U2809 (.Y(n496), 
	.B1(n31), 
	.B0(key_mem[1389]), 
	.A1(n30), 
	.A0(FE_PHN981_key_mem_1261_));
   AOI222X1 U2810 (.Y(n499), 
	.C1(n23), 
	.C0(key_mem[237]), 
	.B1(n22), 
	.B0(key_mem[109]), 
	.A1(n21), 
	.A0(FE_PHN1618_key_mem_365_));
   AOI222X1 U2811 (.Y(n498), 
	.C1(n2800), 
	.C0(key_mem[621]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[493]), 
	.A1(n2823), 
	.A0(FE_PHN1500_key_mem_749_));
   NAND4X1 U2812 (.Y(round_key[4]), 
	.D(n251), 
	.C(n250), 
	.B(n249), 
	.A(n248));
   AOI22X1 U2813 (.Y(n248), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1284]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN775_key_mem_1156_));
   AOI222X1 U2814 (.Y(n251), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[132]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[4]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1738_key_mem_260_));
   AOI222X1 U2815 (.Y(n250), 
	.C1(n2806), 
	.C0(key_mem[516]), 
	.B1(n2818), 
	.B0(key_mem[388]), 
	.A1(n2829), 
	.A0(FE_PHN1809_key_mem_644_));
   NAND4X1 U2816 (.Y(round_key[35]), 
	.D(n315), 
	.C(n314), 
	.B(n313), 
	.A(n312));
   AOI22X1 U2817 (.Y(n312), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1315]), 
	.A1(FE_OFN101_n30), 
	.A0(key_mem[1187]));
   AOI222X1 U2818 (.Y(n315), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[163]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[35]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1735_key_mem_291_));
   AOI222X1 U2819 (.Y(n314), 
	.C1(FE_OFN100_n2800), 
	.C0(key_mem[547]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[419]), 
	.A1(n2827), 
	.A0(FE_PHN1749_key_mem_675_));
   NAND4X1 U2820 (.Y(round_key[107]), 
	.D(n507), 
	.C(n506), 
	.B(n505), 
	.A(n504));
   AOI22X1 U2821 (.Y(n504), 
	.B1(n31), 
	.B0(key_mem[1387]), 
	.A1(n30), 
	.A0(FE_PHN1009_key_mem_1259_));
   AOI222X1 U2822 (.Y(n507), 
	.C1(n23), 
	.C0(key_mem[235]), 
	.B1(n22), 
	.B0(key_mem[107]), 
	.A1(n21), 
	.A0(FE_PHN1677_key_mem_363_));
   AOI222X1 U2823 (.Y(n506), 
	.C1(n2800), 
	.C0(key_mem[619]), 
	.B1(FE_OFN99_n2811), 
	.B0(key_mem[491]), 
	.A1(n2823), 
	.A0(key_mem[747]));
   NAND4X1 U2824 (.Y(round_key[42]), 
	.D(n283), 
	.C(n282), 
	.B(n281), 
	.A(n280));
   AOI22X1 U2825 (.Y(n280), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1322]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN696_key_mem_1194_));
   AOI222X1 U2826 (.Y(n283), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[170]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[42]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1586_key_mem_298_));
   AOI222X1 U2827 (.Y(n282), 
	.C1(n2806), 
	.C0(key_mem[554]), 
	.B1(n2817), 
	.B0(key_mem[426]), 
	.A1(n2828), 
	.A0(FE_PHN1747_key_mem_682_));
   NAND4X1 U2828 (.Y(round_key[65]), 
	.D(n183), 
	.C(n182), 
	.B(n181), 
	.A(n180));
   AOI22X1 U2829 (.Y(n180), 
	.B1(FE_OFN102_n31), 
	.B0(FE_PHN774_key_mem_1345_), 
	.A1(FE_OFN101_n30), 
	.A0(key_mem[1217]));
   AOI222X1 U2830 (.Y(n183), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[193]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[65]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1621_key_mem_321_));
   AOI222X1 U2831 (.Y(n182), 
	.C1(n2800), 
	.C0(key_mem[577]), 
	.B1(n2818), 
	.B0(key_mem[449]), 
	.A1(n2828), 
	.A0(FE_PHN1574_key_mem_705_));
   NAND4X1 U2832 (.Y(round_key[99]), 
	.D(n35), 
	.C(n34), 
	.B(n33), 
	.A(n32));
   AOI22X1 U2833 (.Y(n32), 
	.B1(FE_OFN102_n31), 
	.B0(FE_PHN932_key_mem_1379_), 
	.A1(FE_OFN101_n30), 
	.A0(key_mem[1251]));
   AOI222X1 U2834 (.Y(n35), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[227]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[99]), 
	.A1(n21), 
	.A0(FE_PHN1619_key_mem_355_));
   AOI222X1 U2835 (.Y(n33), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[995]), 
	.B1(n2775), 
	.B0(key_mem[867]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1781_key_mem_1123_));
   NAND4X1 U2836 (.Y(round_key[96]), 
	.D(n47), 
	.C(n46), 
	.B(n45), 
	.A(n44));
   AOI22X1 U2837 (.Y(n44), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1376]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN691_key_mem_1248_));
   AOI222X1 U2838 (.Y(n47), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[224]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[96]), 
	.A1(n21), 
	.A0(FE_PHN1844_key_mem_352_));
   AOI222X1 U2839 (.Y(n45), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[992]), 
	.B1(n2775), 
	.B0(key_mem[864]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1740_key_mem_1120_));
   NAND4X1 U2840 (.Y(round_key[59]), 
	.D(n211), 
	.C(n210), 
	.B(n209), 
	.A(n208));
   AOI22X1 U2841 (.Y(n208), 
	.B1(n31), 
	.B0(key_mem[1339]), 
	.A1(n30), 
	.A0(FE_PHN765_key_mem_1211_));
   AOI222X1 U2842 (.Y(n211), 
	.C1(n23), 
	.C0(key_mem[187]), 
	.B1(n22), 
	.B0(key_mem[59]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1635_key_mem_315_));
   AOI222X1 U2843 (.Y(n209), 
	.C1(n2770), 
	.C0(key_mem[955]), 
	.B1(n2781), 
	.B0(key_mem[827]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1857_key_mem_1083_));
   NAND4X1 U2844 (.Y(round_key[91]), 
	.D(n67), 
	.C(n66), 
	.B(n65), 
	.A(n64));
   AOI22X1 U2845 (.Y(n64), 
	.B1(n31), 
	.B0(key_mem[1371]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN771_key_mem_1243_));
   AOI222X1 U2846 (.Y(n67), 
	.C1(n23), 
	.C0(key_mem[219]), 
	.B1(n22), 
	.B0(key_mem[91]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1572_key_mem_347_));
   AOI222X1 U2847 (.Y(n65), 
	.C1(n2773), 
	.C0(key_mem[987]), 
	.B1(n2775), 
	.B0(key_mem[859]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1823_key_mem_1115_));
   NAND4X1 U2848 (.Y(round_key[27]), 
	.D(n351), 
	.C(n350), 
	.B(n349), 
	.A(n348));
   AOI22X1 U2849 (.Y(n348), 
	.B1(n31), 
	.B0(key_mem[1307]), 
	.A1(n30), 
	.A0(FE_PHN760_key_mem_1179_));
   AOI222X1 U2850 (.Y(n351), 
	.C1(n23), 
	.C0(key_mem[155]), 
	.B1(n22), 
	.B0(key_mem[27]), 
	.A1(n21), 
	.A0(FE_PHN1518_key_mem_283_));
   AOI222X1 U2851 (.Y(n349), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[923]), 
	.B1(n2775), 
	.B0(key_mem[795]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1784_key_mem_1051_));
   NAND4X1 U2852 (.Y(round_key[123]), 
	.D(n435), 
	.C(n434), 
	.B(n433), 
	.A(n432));
   AOI22X1 U2853 (.Y(n432), 
	.B1(n31), 
	.B0(key_mem[1403]), 
	.A1(n30), 
	.A0(key_mem[1275]));
   AOI222X1 U2854 (.Y(n435), 
	.C1(n23), 
	.C0(key_mem[251]), 
	.B1(n22), 
	.B0(key_mem[123]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN755_key_mem_379_));
   AOI222X1 U2855 (.Y(n433), 
	.C1(n2766), 
	.C0(key_mem[1019]), 
	.B1(n2775), 
	.B0(key_mem[891]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1805_key_mem_1147_));
   NAND4X1 U2856 (.Y(round_key[26]), 
	.D(n355), 
	.C(n354), 
	.B(n353), 
	.A(n352));
   AOI22X1 U2857 (.Y(n352), 
	.B1(n31), 
	.B0(key_mem[1306]), 
	.A1(n30), 
	.A0(key_mem[1178]));
   AOI222X1 U2858 (.Y(n355), 
	.C1(n23), 
	.C0(key_mem[154]), 
	.B1(n22), 
	.B0(key_mem[26]), 
	.A1(n21), 
	.A0(FE_PHN1554_key_mem_282_));
   AOI222X1 U2859 (.Y(n353), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[922]), 
	.B1(n2775), 
	.B0(key_mem[794]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1772_key_mem_1050_));
   NAND4X1 U2860 (.Y(round_key[122]), 
	.D(n439), 
	.C(n438), 
	.B(n437), 
	.A(n436));
   AOI22X1 U2861 (.Y(n436), 
	.B1(n31), 
	.B0(key_mem[1402]), 
	.A1(n30), 
	.A0(FE_PHN766_key_mem_1274_));
   AOI222X1 U2862 (.Y(n439), 
	.C1(n23), 
	.C0(key_mem[250]), 
	.B1(n22), 
	.B0(key_mem[122]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1589_key_mem_378_));
   AOI222X1 U2863 (.Y(n437), 
	.C1(n2766), 
	.C0(key_mem[1018]), 
	.B1(n2775), 
	.B0(key_mem[890]), 
	.A1(FE_OFN103_n27), 
	.A0(key_mem[1146]));
   NAND4X1 U2864 (.Y(round_key[90]), 
	.D(n71), 
	.C(n70), 
	.B(n69), 
	.A(n68));
   AOI22X1 U2865 (.Y(n68), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1370]), 
	.A1(n30), 
	.A0(FE_PHN767_key_mem_1242_));
   AOI222X1 U2866 (.Y(n71), 
	.C1(n23), 
	.C0(key_mem[218]), 
	.B1(n22), 
	.B0(key_mem[90]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1690_key_mem_346_));
   AOI222X1 U2867 (.Y(n69), 
	.C1(n2773), 
	.C0(key_mem[986]), 
	.B1(n2775), 
	.B0(key_mem[858]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1885_key_mem_1114_));
   NAND4X1 U2868 (.Y(round_key[58]), 
	.D(n215), 
	.C(n214), 
	.B(n213), 
	.A(n212));
   AOI22X1 U2869 (.Y(n212), 
	.B1(n31), 
	.B0(key_mem[1338]), 
	.A1(n30), 
	.A0(key_mem[1210]));
   AOI222X1 U2870 (.Y(n215), 
	.C1(n23), 
	.C0(key_mem[186]), 
	.B1(n22), 
	.B0(key_mem[58]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1529_key_mem_314_));
   AOI222X1 U2871 (.Y(n213), 
	.C1(n2770), 
	.C0(key_mem[954]), 
	.B1(n2781), 
	.B0(key_mem[826]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1930_key_mem_1082_));
   NAND4X1 U2872 (.Y(round_key[57]), 
	.D(n219), 
	.C(n218), 
	.B(n217), 
	.A(n216));
   AOI22X1 U2873 (.Y(n216), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1337]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN783_key_mem_1209_));
   AOI222X1 U2874 (.Y(n219), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[185]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[57]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1584_key_mem_313_));
   AOI222X1 U2875 (.Y(n217), 
	.C1(n2770), 
	.C0(key_mem[953]), 
	.B1(n2781), 
	.B0(key_mem[825]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1783_key_mem_1081_));
   NAND4X1 U2876 (.Y(round_key[25]), 
	.D(n359), 
	.C(n358), 
	.B(n357), 
	.A(n356));
   AOI22X1 U2877 (.Y(n356), 
	.B1(n31), 
	.B0(FE_PHN2829_key_mem_1305_), 
	.A1(n30), 
	.A0(FE_PHN791_key_mem_1177_));
   AOI222X1 U2878 (.Y(n359), 
	.C1(n23), 
	.C0(key_mem[153]), 
	.B1(n22), 
	.B0(key_mem[25]), 
	.A1(n21), 
	.A0(FE_PHN1623_key_mem_281_));
   AOI222X1 U2879 (.Y(n357), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[921]), 
	.B1(n2775), 
	.B0(key_mem[793]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1876_key_mem_1049_));
   NAND4X1 U2880 (.Y(round_key[121]), 
	.D(n443), 
	.C(n442), 
	.B(n441), 
	.A(n440));
   AOI22X1 U2881 (.Y(n440), 
	.B1(n31), 
	.B0(FE_PHN2834_key_mem_1401_), 
	.A1(n30), 
	.A0(FE_PHN802_key_mem_1273_));
   AOI222X1 U2882 (.Y(n443), 
	.C1(n23), 
	.C0(key_mem[249]), 
	.B1(n22), 
	.B0(key_mem[121]), 
	.A1(n21), 
	.A0(FE_PHN1515_key_mem_377_));
   AOI222X1 U2883 (.Y(n441), 
	.C1(n2766), 
	.C0(key_mem[1017]), 
	.B1(n2775), 
	.B0(FE_PHN3270_key_mem_889_), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1762_key_mem_1145_));
   NAND4X1 U2884 (.Y(round_key[89]), 
	.D(n79), 
	.C(n78), 
	.B(n77), 
	.A(n76));
   AOI22X1 U2885 (.Y(n76), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1369]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN770_key_mem_1241_));
   AOI222X1 U2886 (.Y(n79), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[217]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[89]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1739_key_mem_345_));
   AOI222X1 U2887 (.Y(n77), 
	.C1(n2773), 
	.C0(key_mem[985]), 
	.B1(n2775), 
	.B0(key_mem[857]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1818_key_mem_1113_));
   NAND4X1 U2888 (.Y(round_key[88]), 
	.D(n83), 
	.C(n82), 
	.B(n81), 
	.A(n80));
   AOI22X1 U2889 (.Y(n80), 
	.B1(FE_OFN102_n31), 
	.B0(FE_PHN2830_key_mem_1368_), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN817_key_mem_1240_));
   AOI222X1 U2890 (.Y(n83), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[216]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[88]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1775_key_mem_344_));
   AOI222X1 U2891 (.Y(n81), 
	.C1(n2773), 
	.C0(key_mem[984]), 
	.B1(n2775), 
	.B0(FE_PHN3207_key_mem_856_), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1860_key_mem_1112_));
   NAND4X1 U2892 (.Y(round_key[24]), 
	.D(n363), 
	.C(n362), 
	.B(n361), 
	.A(n360));
   AOI22X1 U2893 (.Y(n360), 
	.B1(n31), 
	.B0(FE_PHN2827_key_mem_1304_), 
	.A1(n30), 
	.A0(FE_PHN819_key_mem_1176_));
   AOI222X1 U2894 (.Y(n363), 
	.C1(n23), 
	.C0(key_mem[152]), 
	.B1(n22), 
	.B0(key_mem[24]), 
	.A1(n21), 
	.A0(FE_PHN1634_key_mem_280_));
   AOI222X1 U2895 (.Y(n361), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[920]), 
	.B1(n2775), 
	.B0(key_mem[792]), 
	.A1(FE_OFN103_n27), 
	.A0(key_mem[1048]));
   NAND4X1 U2896 (.Y(round_key[120]), 
	.D(n447), 
	.C(n446), 
	.B(n445), 
	.A(n444));
   AOI22X1 U2897 (.Y(n444), 
	.B1(n31), 
	.B0(FE_PHN3229_key_mem_1400_), 
	.A1(n30), 
	.A0(FE_PHN1899_key_mem_1272_));
   AOI222X1 U2898 (.Y(n447), 
	.C1(n23), 
	.C0(key_mem[248]), 
	.B1(n22), 
	.B0(key_mem[120]), 
	.A1(n21), 
	.A0(FE_PHN1849_key_mem_376_));
   AOI222X1 U2899 (.Y(n445), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[1016]), 
	.B1(n2775), 
	.B0(key_mem[888]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1858_key_mem_1144_));
   NAND4X1 U2900 (.Y(round_key[127]), 
	.D(n419), 
	.C(n418), 
	.B(n417), 
	.A(n416));
   AOI22X1 U2901 (.Y(n416), 
	.B1(n31), 
	.B0(FE_PHN3444_key_mem_1407_), 
	.A1(n30), 
	.A0(FE_PHN3091_key_mem_1279_));
   AOI222X1 U2902 (.Y(n419), 
	.C1(n23), 
	.C0(FE_PHN3418_key_mem_255_), 
	.B1(n22), 
	.B0(FE_PHN3208_key_mem_127_), 
	.A1(n21), 
	.A0(FE_PHN1517_key_mem_383_));
   AOI222X1 U2903 (.Y(n417), 
	.C1(n2766), 
	.C0(key_mem[1023]), 
	.B1(n2775), 
	.B0(FE_PHN3275_key_mem_895_), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1884_key_mem_1151_));
   NAND4X1 U2904 (.Y(round_key[126]), 
	.D(n423), 
	.C(n422), 
	.B(n421), 
	.A(n420));
   AOI22X1 U2905 (.Y(n420), 
	.B1(n31), 
	.B0(key_mem[1406]), 
	.A1(n30), 
	.A0(FE_PHN1766_key_mem_1278_));
   AOI222X1 U2906 (.Y(n423), 
	.C1(n23), 
	.C0(key_mem[254]), 
	.B1(n22), 
	.B0(FE_PHN3089_key_mem_126_), 
	.A1(n21), 
	.A0(FE_PHN1503_key_mem_382_));
   AOI222X1 U2907 (.Y(n421), 
	.C1(n2766), 
	.C0(key_mem[1022]), 
	.B1(n2775), 
	.B0(key_mem[894]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1814_key_mem_1150_));
   NAND4X1 U2908 (.Y(round_key[125]), 
	.D(n427), 
	.C(n426), 
	.B(n425), 
	.A(n424));
   AOI22X1 U2909 (.Y(n424), 
	.B1(n31), 
	.B0(key_mem[1405]), 
	.A1(n30), 
	.A0(FE_PHN792_key_mem_1277_));
   AOI222X1 U2910 (.Y(n427), 
	.C1(n23), 
	.C0(key_mem[253]), 
	.B1(n22), 
	.B0(key_mem[125]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1501_key_mem_381_));
   AOI222X1 U2911 (.Y(n425), 
	.C1(n2766), 
	.C0(key_mem[1021]), 
	.B1(n2775), 
	.B0(key_mem[893]), 
	.A1(FE_OFN103_n27), 
	.A0(key_mem[1149]));
   NAND4X1 U2912 (.Y(round_key[92]), 
	.D(n63), 
	.C(n62), 
	.B(n61), 
	.A(n60));
   AOI22X1 U2913 (.Y(n60), 
	.B1(FE_OFN102_n31), 
	.B0(FE_PHN788_key_mem_1372_), 
	.A1(FE_OFN101_n30), 
	.A0(key_mem[1244]));
   AOI222X1 U2914 (.Y(n63), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[220]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[92]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1725_key_mem_348_));
   AOI222X1 U2915 (.Y(n61), 
	.C1(n2773), 
	.C0(key_mem[988]), 
	.B1(n2775), 
	.B0(key_mem[860]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1843_key_mem_1116_));
   NAND4X1 U2916 (.Y(round_key[56]), 
	.D(n223), 
	.C(n222), 
	.B(n221), 
	.A(n220));
   AOI22X1 U2917 (.Y(n220), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1336]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN786_key_mem_1208_));
   AOI222X1 U2918 (.Y(n223), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[184]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[56]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1537_key_mem_312_));
   AOI222X1 U2919 (.Y(n221), 
	.C1(n2770), 
	.C0(key_mem[952]), 
	.B1(n2781), 
	.B0(key_mem[824]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1730_key_mem_1080_));
   NAND4X1 U2920 (.Y(round_key[63]), 
	.D(n191), 
	.C(n190), 
	.B(n189), 
	.A(n188));
   AOI22X1 U2921 (.Y(n188), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1343]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN1700_key_mem_1215_));
   AOI222X1 U2922 (.Y(n191), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[191]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[63]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1496_key_mem_319_));
   AOI222X1 U2923 (.Y(n189), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[959]), 
	.B1(n2781), 
	.B0(key_mem[831]), 
	.A1(FE_OFN104_n27), 
	.A0(key_mem[1087]));
   NAND4X1 U2924 (.Y(round_key[62]), 
	.D(n195), 
	.C(n194), 
	.B(n193), 
	.A(n192));
   AOI22X1 U2925 (.Y(n192), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1342]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN800_key_mem_1214_));
   AOI222X1 U2926 (.Y(n195), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[190]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[62]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1806_key_mem_318_));
   AOI222X1 U2927 (.Y(n193), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[958]), 
	.B1(n2781), 
	.B0(key_mem[830]), 
	.A1(FE_OFN104_n27), 
	.A0(key_mem[1086]));
   NAND4X1 U2928 (.Y(round_key[61]), 
	.D(n199), 
	.C(n198), 
	.B(n197), 
	.A(n196));
   AOI22X1 U2929 (.Y(n196), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1341]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN782_key_mem_1213_));
   AOI222X1 U2930 (.Y(n199), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[189]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[61]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1658_key_mem_317_));
   AOI222X1 U2931 (.Y(n197), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[957]), 
	.B1(n2781), 
	.B0(key_mem[829]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1856_key_mem_1085_));
   NAND4X1 U2932 (.Y(round_key[60]), 
	.D(n203), 
	.C(n202), 
	.B(n201), 
	.A(n200));
   AOI22X1 U2933 (.Y(n200), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1340]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN797_key_mem_1212_));
   AOI222X1 U2934 (.Y(n203), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[188]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[60]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1710_key_mem_316_));
   AOI222X1 U2935 (.Y(n201), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[956]), 
	.B1(n2781), 
	.B0(key_mem[828]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1835_key_mem_1084_));
   NAND4X1 U2936 (.Y(round_key[28]), 
	.D(n347), 
	.C(n346), 
	.B(n345), 
	.A(n344));
   AOI22X1 U2937 (.Y(n344), 
	.B1(n31), 
	.B0(key_mem[1308]), 
	.A1(n30), 
	.A0(key_mem[1180]));
   AOI222X1 U2938 (.Y(n347), 
	.C1(n23), 
	.C0(key_mem[156]), 
	.B1(n22), 
	.B0(key_mem[28]), 
	.A1(n21), 
	.A0(FE_PHN1482_key_mem_284_));
   AOI222X1 U2939 (.Y(n345), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[924]), 
	.B1(n2780), 
	.B0(key_mem[796]), 
	.A1(FE_OFN103_n27), 
	.A0(key_mem[1052]));
   NAND4X1 U2940 (.Y(round_key[124]), 
	.D(n431), 
	.C(n430), 
	.B(n429), 
	.A(n428));
   AOI22X1 U2941 (.Y(n428), 
	.B1(n31), 
	.B0(key_mem[1404]), 
	.A1(n30), 
	.A0(FE_PHN780_key_mem_1276_));
   AOI222X1 U2942 (.Y(n431), 
	.C1(n23), 
	.C0(key_mem[252]), 
	.B1(n22), 
	.B0(key_mem[124]), 
	.A1(FE_OFN108_n21), 
	.A0(FE_PHN1670_key_mem_380_));
   AOI222X1 U2943 (.Y(n429), 
	.C1(n2766), 
	.C0(key_mem[1020]), 
	.B1(n2775), 
	.B0(key_mem[892]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1808_key_mem_1148_));
   NAND4X1 U2944 (.Y(round_key[31]), 
	.D(n331), 
	.C(n330), 
	.B(n329), 
	.A(n328));
   AOI22X1 U2945 (.Y(n328), 
	.B1(n31), 
	.B0(FE_PHN1834_key_mem_1311_), 
	.A1(n30), 
	.A0(FE_PHN3319_key_mem_1183_));
   AOI222X1 U2946 (.Y(n331), 
	.C1(n23), 
	.C0(FE_PHN3411_key_mem_159_), 
	.B1(n22), 
	.B0(FE_PHN3085_key_mem_31_), 
	.A1(n21), 
	.A0(FE_PHN764_key_mem_287_));
   AOI222X1 U2947 (.Y(n329), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[927]), 
	.B1(n2780), 
	.B0(FE_PHN3210_key_mem_799_), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1864_key_mem_1055_));
   NAND4X1 U2948 (.Y(round_key[30]), 
	.D(n335), 
	.C(n334), 
	.B(n333), 
	.A(n332));
   AOI22X1 U2949 (.Y(n332), 
	.B1(n31), 
	.B0(key_mem[1310]), 
	.A1(n30), 
	.A0(FE_PHN808_key_mem_1182_));
   AOI222X1 U2950 (.Y(n335), 
	.C1(n23), 
	.C0(key_mem[158]), 
	.B1(n22), 
	.B0(key_mem[30]), 
	.A1(n21), 
	.A0(FE_PHN1477_key_mem_286_));
   AOI222X1 U2951 (.Y(n333), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[926]), 
	.B1(n2780), 
	.B0(key_mem[798]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1769_key_mem_1054_));
   NAND4X1 U2952 (.Y(round_key[29]), 
	.D(n343), 
	.C(n342), 
	.B(n341), 
	.A(n340));
   AOI22X1 U2953 (.Y(n340), 
	.B1(n31), 
	.B0(key_mem[1309]), 
	.A1(n30), 
	.A0(key_mem[1181]));
   AOI222X1 U2954 (.Y(n343), 
	.C1(n23), 
	.C0(key_mem[157]), 
	.B1(n22), 
	.B0(key_mem[29]), 
	.A1(n21), 
	.A0(FE_PHN1802_key_mem_285_));
   AOI222X1 U2955 (.Y(n341), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[925]), 
	.B1(n2780), 
	.B0(key_mem[797]), 
	.A1(FE_OFN103_n27), 
	.A0(FE_PHN1868_key_mem_1053_));
   NAND4X1 U2956 (.Y(round_key[94]), 
	.D(n55), 
	.C(n54), 
	.B(n53), 
	.A(n52));
   AOI22X1 U2957 (.Y(n52), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1374]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN794_key_mem_1246_));
   AOI222X1 U2958 (.Y(n55), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[222]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[94]), 
	.A1(n21), 
	.A0(FE_PHN1614_key_mem_350_));
   AOI222X1 U2959 (.Y(n53), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[990]), 
	.B1(n2775), 
	.B0(key_mem[862]), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1803_key_mem_1118_));
   NAND4X1 U2960 (.Y(round_key[93]), 
	.D(n59), 
	.C(n58), 
	.B(n57), 
	.A(n56));
   AOI22X1 U2961 (.Y(n56), 
	.B1(FE_OFN102_n31), 
	.B0(key_mem[1373]), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN773_key_mem_1245_));
   AOI222X1 U2962 (.Y(n59), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[221]), 
	.B1(FE_OFN106_n22), 
	.B0(key_mem[93]), 
	.A1(FE_OFN107_n21), 
	.A0(FE_PHN1851_key_mem_349_));
   AOI222X1 U2963 (.Y(n57), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[989]), 
	.B1(n2775), 
	.B0(key_mem[861]), 
	.A1(FE_OFN103_n27), 
	.A0(key_mem[1117]));
   NAND4X1 U2964 (.Y(round_key[95]), 
	.D(n51), 
	.C(n50), 
	.B(n49), 
	.A(n48));
   AOI22X1 U2965 (.Y(n48), 
	.B1(FE_OFN102_n31), 
	.B0(FE_PHN2833_key_mem_1375_), 
	.A1(FE_OFN101_n30), 
	.A0(FE_PHN811_key_mem_1247_));
   AOI222X1 U2966 (.Y(n51), 
	.C1(FE_OFN109_n23), 
	.C0(key_mem[223]), 
	.B1(FE_OFN106_n22), 
	.B0(FE_PHN3201_key_mem_95_), 
	.A1(n21), 
	.A0(FE_PHN1754_key_mem_351_));
   AOI222X1 U2967 (.Y(n49), 
	.C1(FE_OFN105_n2763), 
	.C0(key_mem[991]), 
	.B1(n2775), 
	.B0(FE_PHN3203_key_mem_863_), 
	.A1(FE_OFN104_n27), 
	.A0(FE_PHN1817_key_mem_1119_));
   NOR4BX1 U2969 (.Y(n27), 
	.D(round[3]), 
	.C(round[2]), 
	.B(n2877), 
	.AN(n2876));
   OR3XL U2970 (.Y(n4), 
	.C(n2876), 
	.B(round[2]), 
	.A(n2877));
   OR3XL U2971 (.Y(n5), 
	.C(n2878), 
	.B(round[1]), 
	.A(round[0]));
   OR3XL U2972 (.Y(n7), 
	.C(n2878), 
	.B(round[1]), 
	.A(n2876));
   OR3XL U2973 (.Y(n8), 
	.C(n2878), 
	.B(round[0]), 
	.A(n2877));
   NOR2BX4 U2974 (.Y(n31), 
	.B(round[0]), 
	.AN(n540));
   NOR3X1 U2975 (.Y(n673), 
	.C(n675), 
	.B(FE_PHN116_round_ctr_reg_3_), 
	.A(FE_PHN178_round_ctr_reg_2_));
   NAND3X1 U2976 (.Y(n672), 
	.C(FE_PHN198_round_ctr_reg_0_), 
	.B(n2872), 
	.A(n673));
   NAND3X1 U2977 (.Y(n674), 
	.C(FE_PHN112_round_ctr_reg_1_), 
	.B(FE_PHN411_n6), 
	.A(n673));
   OAI221XL U2978 (.Y(n884), 
	.C0(n2870), 
	.B1(n2879), 
	.B0(FE_PHN120_key_mem_ctrl_reg_1_), 
	.A1(FE_PHN254_n689), 
	.A0(n2871));
   INVX1 U2979 (.Y(n2879), 
	.A(init));
   OAI32XL U2980 (.Y(n2423), 
	.B1(n2872), 
	.B0(n2869), 
	.A2(n675), 
	.A1(FE_PHN112_round_ctr_reg_1_), 
	.A0(FE_PHN411_n6));
   INVX1 U2981 (.Y(n2871), 
	.A(FE_PHN120_key_mem_ctrl_reg_1_));
   XOR2X1 U2982 (.Y(n765), 
	.B(FE_PHN940_prev_key1_reg_95_), 
	.A(FE_PHN1434_prev_key1_reg_127_));
   XOR2X1 U2983 (.Y(n786), 
	.B(FE_PHN979_prev_key1_reg_88_), 
	.A(FE_PHN1416_prev_key1_reg_120_));
   XOR2X1 U2984 (.Y(n768), 
	.B(FE_PHN933_prev_key1_reg_94_), 
	.A(prev_key1_reg[126]));
   XOR2X1 U2985 (.Y(n771), 
	.B(FE_PHN757_prev_key1_reg_93_), 
	.A(FE_PHN1391_prev_key1_reg_125_));
   XOR2X1 U2986 (.Y(n774), 
	.B(FE_PHN919_prev_key1_reg_92_), 
	.A(FE_PHN1421_prev_key1_reg_124_));
   XOR2X1 U2987 (.Y(n777), 
	.B(FE_PHN921_prev_key1_reg_91_), 
	.A(FE_PHN1413_prev_key1_reg_123_));
   XOR2X1 U2988 (.Y(n780), 
	.B(FE_PHN924_prev_key1_reg_90_), 
	.A(FE_PHN1392_prev_key1_reg_122_));
   XOR2X1 U2989 (.Y(n783), 
	.B(FE_PHN922_prev_key1_reg_89_), 
	.A(FE_PHN1395_prev_key1_reg_121_));
   NAND2X1 U2990 (.Y(n880), 
	.B(FE_PHN290_key_mem_ctrl_reg_0_), 
	.A(n2871));
   INVX1 U2991 (.Y(n2869), 
	.A(n878));
   OAI21XL U2992 (.Y(n878), 
	.B0(n879), 
	.A1(n675), 
	.A0(FE_PHN198_round_ctr_reg_0_));
   OAI2BB1X1 U2993 (.Y(n2422), 
	.B0(n877), 
	.A1N(FE_PHN178_round_ctr_reg_2_), 
	.A0N(n876));
   NAND4XL U2994 (.Y(n877), 
	.D(n2873), 
	.C(FE_PHN155_n3), 
	.B(FE_PHN198_round_ctr_reg_0_), 
	.A(FE_PHN112_round_ctr_reg_1_));
   NAND2BX1 U2995 (.Y(n2431), 
	.B(FE_PHN155_n3), 
	.AN(FE_PHN1989_rcon_reg_6_));
   NAND2BX1 U2996 (.Y(n2428), 
	.B(FE_PHN155_n3), 
	.AN(FE_PHN1263_rcon_reg_1_));
   NAND2X1 U2997 (.Y(n2427), 
	.B(FE_PHN155_n3), 
	.A(n882));
   XOR2X1 U2998 (.Y(n882), 
	.B(n2875), 
	.A(FE_PHN1033_rcon_reg_2_));
   AND2X2 U2999 (.Y(n2424), 
	.B(FE_PHN155_n3), 
	.A(FE_PHN1241_rcon_reg_5_));
   AND2X2 U3000 (.Y(n2425), 
	.B(FE_PHN155_n3), 
	.A(FE_PHN1257_rcon_reg_4_));
   INVX1 U3001 (.Y(n2875), 
	.A(FE_PHN912_rcon_reg_7_));
   NAND3X1 U3002 (.Y(n542), 
	.C(init), 
	.B(n2871), 
	.A(n2870));
   NOR2X1 U3003 (.Y(n2426), 
	.B(n675), 
	.A(FE_PHN3406_n881));
   XOR2X1 U3004 (.Y(n881), 
	.B(n2875), 
	.A(FE_PHN1036_rcon_reg_3_));
   NOR2X1 U3005 (.Y(n2429), 
	.B(n675), 
	.A(FE_PHN3407_n883));
   XOR2X1 U3006 (.Y(n883), 
	.B(n2875), 
	.A(FE_PHN1034_rcon_reg_0_));
   INVX1 U3007 (.Y(n2868), 
	.A(n541));
   AOI22X1 U3008 (.Y(n541), 
	.B1(ready), 
	.B0(n542), 
	.A1(FE_PHN290_key_mem_ctrl_reg_0_), 
	.A0(FE_PHN120_key_mem_ctrl_reg_1_));
endmodule

module aes_sbox (
	sboxw, 
	new_sboxw);
   input [31:0] sboxw;
   output [31:0] new_sboxw;

   // Internal wires
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n227;
   wire n228;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n242;
   wire n243;
   wire n244;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n274;
   wire n275;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire n556;
   wire n557;
   wire n558;
   wire n559;
   wire n560;
   wire n561;
   wire n562;
   wire n563;
   wire n564;
   wire n565;
   wire n566;
   wire n567;
   wire n568;
   wire n569;
   wire n570;
   wire n572;
   wire n573;
   wire n574;
   wire n575;
   wire n576;
   wire n577;
   wire n578;
   wire n579;
   wire n580;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire n593;
   wire n594;
   wire n595;
   wire n596;
   wire n597;
   wire n598;
   wire n599;
   wire n600;
   wire n601;
   wire n602;
   wire n603;
   wire n604;
   wire n605;
   wire n606;
   wire n607;
   wire n608;
   wire n609;
   wire n610;
   wire n611;
   wire n612;
   wire n613;
   wire n614;
   wire n615;
   wire n616;
   wire n617;
   wire n618;
   wire n619;
   wire n620;
   wire n621;
   wire n622;
   wire n623;
   wire n624;
   wire n625;
   wire n626;
   wire n627;
   wire n628;
   wire n629;
   wire n631;
   wire n632;
   wire n633;
   wire n634;
   wire n636;
   wire n637;
   wire n638;
   wire n639;
   wire n640;
   wire n641;
   wire n642;
   wire n643;
   wire n644;
   wire n646;
   wire n647;
   wire n648;
   wire n649;
   wire n650;
   wire n651;
   wire n652;
   wire n653;
   wire n654;
   wire n655;
   wire n656;
   wire n657;
   wire n658;
   wire n659;
   wire n660;
   wire n661;
   wire n662;
   wire n663;
   wire n664;
   wire n665;
   wire n666;
   wire n667;
   wire n668;
   wire n669;
   wire n670;
   wire n671;
   wire n673;
   wire n674;
   wire n675;
   wire n676;
   wire n677;
   wire n678;
   wire n679;
   wire n680;
   wire n681;
   wire n682;
   wire n683;
   wire n684;
   wire n685;
   wire n686;
   wire n687;
   wire n688;
   wire n689;
   wire n690;
   wire n691;
   wire n692;
   wire n693;
   wire n694;
   wire n695;
   wire n696;
   wire n697;
   wire n698;
   wire n699;
   wire n700;
   wire n701;
   wire n702;
   wire n703;
   wire n704;
   wire n705;
   wire n706;
   wire n707;
   wire n708;
   wire n709;
   wire n710;
   wire n711;
   wire n712;
   wire n713;
   wire n714;
   wire n715;
   wire n716;
   wire n717;
   wire n718;
   wire n719;
   wire n720;
   wire n721;
   wire n722;
   wire n723;
   wire n724;
   wire n725;
   wire n726;
   wire n727;
   wire n728;
   wire n729;
   wire n730;
   wire n731;
   wire n732;
   wire n733;
   wire n734;
   wire n735;
   wire n736;
   wire n737;
   wire n738;
   wire n740;
   wire n741;
   wire n742;
   wire n743;
   wire n744;
   wire n745;
   wire n746;
   wire n747;
   wire n748;
   wire n749;
   wire n750;
   wire n751;
   wire n752;
   wire n753;
   wire n754;
   wire n755;
   wire n756;
   wire n757;
   wire n758;
   wire n759;
   wire n760;
   wire n761;
   wire n762;
   wire n763;
   wire n764;
   wire n765;
   wire n766;
   wire n767;
   wire n768;
   wire n769;
   wire n770;
   wire n771;
   wire n772;
   wire n773;
   wire n774;
   wire n775;
   wire n776;
   wire n777;
   wire n778;
   wire n779;
   wire n780;
   wire n781;
   wire n782;
   wire n783;
   wire n784;
   wire n785;
   wire n786;
   wire n787;
   wire n788;
   wire n789;
   wire n790;
   wire n791;
   wire n792;
   wire n793;
   wire n794;
   wire n795;
   wire n796;
   wire n797;
   wire n798;
   wire n799;
   wire n800;
   wire n801;
   wire n802;
   wire n803;
   wire n804;
   wire n805;
   wire n806;
   wire n807;
   wire n808;
   wire n809;
   wire n810;
   wire n811;
   wire n812;
   wire n813;
   wire n814;
   wire n815;
   wire n816;
   wire n817;
   wire n818;
   wire n819;
   wire n820;
   wire n821;
   wire n822;
   wire n823;
   wire n824;
   wire n825;
   wire n826;
   wire n827;
   wire n828;
   wire n829;
   wire n830;
   wire n831;
   wire n832;
   wire n833;
   wire n834;
   wire n835;
   wire n836;
   wire n837;
   wire n838;
   wire n839;
   wire n840;
   wire n841;
   wire n842;
   wire n843;
   wire n844;
   wire n845;
   wire n846;
   wire n847;
   wire n848;
   wire n849;
   wire n850;
   wire n851;
   wire n852;
   wire n853;
   wire n854;
   wire n855;
   wire n856;
   wire n857;
   wire n858;
   wire n859;
   wire n860;
   wire n861;
   wire n862;
   wire n863;
   wire n864;
   wire n865;
   wire n866;
   wire n867;
   wire n868;
   wire n869;
   wire n870;
   wire n871;
   wire n872;
   wire n873;
   wire n874;
   wire n875;
   wire n876;
   wire n877;
   wire n878;
   wire n879;
   wire n880;
   wire n881;
   wire n882;
   wire n883;
   wire n884;
   wire n885;
   wire n886;
   wire n887;
   wire n888;
   wire n889;
   wire n890;
   wire n891;
   wire n892;
   wire n893;
   wire n894;
   wire n895;
   wire n896;
   wire n897;
   wire n898;
   wire n899;
   wire n900;
   wire n901;
   wire n903;
   wire n904;
   wire n905;
   wire n906;
   wire n907;
   wire n908;
   wire n909;
   wire n910;
   wire n911;
   wire n912;
   wire n913;
   wire n914;
   wire n915;
   wire n916;
   wire n917;
   wire n918;
   wire n919;
   wire n920;
   wire n921;
   wire n922;
   wire n923;
   wire n924;
   wire n926;
   wire n927;
   wire n928;
   wire n929;
   wire n930;
   wire n931;
   wire n932;
   wire n933;
   wire n934;
   wire n935;
   wire n936;
   wire n937;
   wire n938;
   wire n939;
   wire n941;
   wire n942;
   wire n943;
   wire n944;
   wire n945;
   wire n946;
   wire n947;
   wire n948;
   wire n949;
   wire n950;
   wire n951;
   wire n952;
   wire n953;
   wire n954;
   wire n955;
   wire n956;
   wire n957;
   wire n958;
   wire n959;
   wire n960;
   wire n961;
   wire n962;
   wire n963;
   wire n964;
   wire n965;
   wire n966;
   wire n967;
   wire n968;
   wire n969;
   wire n970;
   wire n971;
   wire n972;
   wire n973;
   wire n974;
   wire n975;
   wire n976;
   wire n977;
   wire n978;
   wire n979;
   wire n980;
   wire n981;
   wire n982;
   wire n983;
   wire n985;
   wire n986;
   wire n987;
   wire n988;
   wire n990;
   wire n991;
   wire n992;
   wire n993;
   wire n994;
   wire n995;
   wire n996;
   wire n997;
   wire n998;
   wire n999;
   wire n1000;
   wire n1001;
   wire n1002;
   wire n1003;
   wire n1004;
   wire n1005;
   wire n1006;
   wire n1007;
   wire n1008;
   wire n1009;
   wire n1010;
   wire n1011;
   wire n1012;
   wire n1013;
   wire n1014;
   wire n1015;
   wire n1016;
   wire n1017;
   wire n1018;
   wire n1019;
   wire n1020;
   wire n1021;
   wire n1022;
   wire n1023;
   wire n1024;
   wire n1025;
   wire n1026;
   wire n1027;
   wire n1028;
   wire n1029;
   wire n1030;
   wire n1031;
   wire n1032;
   wire n1033;
   wire n1034;
   wire n1035;
   wire n1036;
   wire n1037;
   wire n1038;
   wire n1039;
   wire n1040;
   wire n1041;
   wire n1042;
   wire n1043;
   wire n1044;
   wire n1045;
   wire n1046;
   wire n1047;
   wire n1048;
   wire n1049;
   wire n1050;
   wire n1051;
   wire n1052;
   wire n1053;
   wire n1054;
   wire n1055;
   wire n1056;
   wire n1057;
   wire n1058;
   wire n1059;
   wire n1062;
   wire n1063;
   wire n1064;
   wire n1065;
   wire n1066;
   wire n1067;
   wire n1068;
   wire n1069;
   wire n1070;
   wire n1071;
   wire n1072;
   wire n1073;
   wire n1074;
   wire n1075;
   wire n1076;
   wire n1077;
   wire n1078;
   wire n1079;
   wire n1080;
   wire n1081;
   wire n1082;
   wire n1083;
   wire n1084;
   wire n1085;
   wire n1086;
   wire n1087;
   wire n1088;
   wire n1089;
   wire n1090;
   wire n1091;
   wire n1092;
   wire n1093;
   wire n1094;
   wire n1095;
   wire n1096;
   wire n1097;
   wire n1098;
   wire n1099;
   wire n1100;
   wire n1101;
   wire n1103;
   wire n1104;
   wire n1105;
   wire n1106;
   wire n1107;
   wire n1108;
   wire n1109;
   wire n1110;
   wire n1111;
   wire n1112;
   wire n1113;
   wire n1114;
   wire n1115;
   wire n1116;
   wire n1117;
   wire n1118;
   wire n1119;
   wire n1120;
   wire n1121;
   wire n1122;
   wire n1123;
   wire n1124;
   wire n1125;
   wire n1126;
   wire n1127;
   wire n1128;
   wire n1129;
   wire n1130;
   wire n1131;
   wire n1132;
   wire n1133;
   wire n1134;
   wire n1135;
   wire n1136;
   wire n1137;
   wire n1138;
   wire n1139;
   wire n1140;
   wire n1141;
   wire n1142;
   wire n1143;
   wire n1144;
   wire n1145;
   wire n1146;
   wire n1147;
   wire n1148;
   wire n1149;
   wire n1150;
   wire n1151;
   wire n1152;
   wire n1153;
   wire n1154;
   wire n1155;
   wire n1156;
   wire n1157;
   wire n1158;
   wire n1159;
   wire n1160;
   wire n1161;
   wire n1162;
   wire n1163;
   wire n1164;
   wire n1165;
   wire n1166;
   wire n1167;
   wire n1168;
   wire n1169;
   wire n1170;
   wire n1171;
   wire n1172;
   wire n1173;
   wire n1174;
   wire n1175;
   wire n1176;
   wire n1177;
   wire n1178;
   wire n1179;
   wire n1180;
   wire n1181;
   wire n1182;
   wire n1183;
   wire n1184;
   wire n1185;
   wire n1186;
   wire n1187;
   wire n1188;
   wire n1189;
   wire n1190;
   wire n1191;
   wire n1192;
   wire n1193;
   wire n1194;
   wire n1195;
   wire n1196;
   wire n1197;
   wire n1198;
   wire n1199;
   wire n1200;
   wire n1201;
   wire n1202;
   wire n1203;
   wire n1204;
   wire n1205;
   wire n1206;
   wire n1207;
   wire n1208;
   wire n1209;
   wire n1210;
   wire n1211;
   wire n1212;
   wire n1213;
   wire n1214;
   wire n1215;
   wire n1216;
   wire n1217;
   wire n1218;
   wire n1219;
   wire n1220;
   wire n1221;
   wire n1222;
   wire n1223;
   wire n1224;
   wire n1225;
   wire n1226;
   wire n1227;
   wire n1228;
   wire n1229;
   wire n1230;
   wire n1231;
   wire n1232;
   wire n1233;
   wire n1234;
   wire n1235;
   wire n1236;
   wire n1237;
   wire n1238;
   wire n1239;
   wire n1240;
   wire n1241;
   wire n1242;
   wire n1243;
   wire n1244;
   wire n1245;
   wire n1246;
   wire n1247;
   wire n1248;
   wire n1249;
   wire n1250;
   wire n1252;
   wire n1253;
   wire n1254;
   wire n1255;
   wire n1256;
   wire n1257;
   wire n1258;
   wire n1259;
   wire n1260;
   wire n1261;
   wire n1262;
   wire n1263;
   wire n1264;
   wire n1265;
   wire n1266;
   wire n1267;
   wire n1268;
   wire n1269;
   wire n1270;
   wire n1271;
   wire n1272;
   wire n1273;
   wire n1274;
   wire n1275;
   wire n1276;
   wire n1277;
   wire n1278;
   wire n1279;
   wire n1280;
   wire n1281;
   wire n1282;
   wire n1283;
   wire n1284;
   wire n1285;
   wire n1286;
   wire n1287;
   wire n1288;
   wire n1289;
   wire n1290;
   wire n1291;
   wire n1292;
   wire n1293;
   wire n1294;
   wire n1295;
   wire n1296;
   wire n1297;
   wire n1298;
   wire n1299;
   wire n1300;
   wire n1301;
   wire n1302;
   wire n1303;
   wire n1304;
   wire n1305;
   wire n1306;
   wire n1307;
   wire n1308;
   wire n1309;
   wire n1310;
   wire n1311;
   wire n1312;
   wire n1313;
   wire n1314;
   wire n1315;
   wire n1316;
   wire n1317;
   wire n1318;
   wire n1319;
   wire n1320;
   wire n1321;
   wire n1322;
   wire n1323;
   wire n1324;
   wire n1325;
   wire n1326;
   wire n1327;
   wire n1328;
   wire n1329;
   wire n1330;
   wire n1331;
   wire n1332;
   wire n1333;
   wire n1334;
   wire n1335;
   wire n1336;
   wire n1337;
   wire n1338;
   wire n1339;
   wire n1340;
   wire n1341;
   wire n1342;
   wire n1343;
   wire n1344;
   wire n1345;
   wire n1346;
   wire n1347;
   wire n1348;
   wire n1349;
   wire n1350;
   wire n1351;
   wire n1352;
   wire n1353;
   wire n1354;
   wire n1355;
   wire n1356;
   wire n1357;
   wire n1358;
   wire n1359;
   wire n1360;
   wire n1361;
   wire n1362;
   wire n1363;
   wire n1364;
   wire n1365;
   wire n1366;
   wire n1367;
   wire n1368;
   wire n1369;
   wire n1370;
   wire n1371;
   wire n1372;
   wire n1373;
   wire n1374;
   wire n1375;
   wire n1376;
   wire n1377;
   wire n1378;
   wire n1379;
   wire n1380;
   wire n1381;
   wire n1382;
   wire n1383;
   wire n1384;
   wire n1385;
   wire n1386;
   wire n1387;
   wire n1388;
   wire n1389;
   wire n1390;
   wire n1391;
   wire n1392;
   wire n1393;
   wire n1394;
   wire n1395;
   wire n1396;
   wire n1397;
   wire n1398;
   wire n1399;
   wire n1400;
   wire n1401;
   wire n1402;
   wire n1403;
   wire n1404;
   wire n1405;
   wire n1406;
   wire n1407;
   wire n1408;
   wire n1409;
   wire n1410;
   wire n1411;
   wire n1412;
   wire n1413;
   wire n1414;
   wire n1415;
   wire n1416;
   wire n1417;
   wire n1418;
   wire n1419;
   wire n1420;
   wire n1421;
   wire n1422;
   wire n1423;
   wire n1424;
   wire n1425;
   wire n1426;
   wire n1427;
   wire n1428;
   wire n1429;
   wire n1430;
   wire n1431;
   wire n1432;
   wire n1433;
   wire n1434;
   wire n1435;
   wire n1436;
   wire n1437;
   wire n1438;
   wire n1439;
   wire n1440;
   wire n1441;
   wire n1442;
   wire n1443;
   wire n1444;
   wire n1445;
   wire n1446;
   wire n1447;
   wire n1448;
   wire n1449;
   wire n1450;
   wire n1451;
   wire n1452;
   wire n1453;
   wire n1454;
   wire n1455;
   wire n1456;
   wire n1457;
   wire n1458;
   wire n1459;
   wire n1460;
   wire n1461;
   wire n1462;
   wire n1463;
   wire n1464;
   wire n1465;
   wire n1466;
   wire n1467;
   wire n1468;
   wire n1469;
   wire n1470;
   wire n1471;
   wire n1472;
   wire n1473;
   wire n1474;
   wire n1475;
   wire n1476;
   wire n1477;
   wire n1478;
   wire n1479;
   wire n1480;
   wire n1481;
   wire n1482;
   wire n1483;
   wire n1484;
   wire n1485;
   wire n1486;
   wire n1487;
   wire n1488;
   wire n1489;
   wire n1490;
   wire n1491;
   wire n1492;
   wire n1493;
   wire n1494;
   wire n1496;
   wire n1497;
   wire n1498;
   wire n1499;
   wire n1500;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n142;
   wire n143;
   wire n146;
   wire n147;
   wire n148;
   wire n150;
   wire n151;
   wire n153;
   wire n156;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n229;
   wire n273;
   wire n276;
   wire n342;
   wire n401;
   wire n406;
   wire n413;
   wire n477;
   wire n478;
   wire n519;
   wire n571;
   wire n630;
   wire n635;
   wire n645;
   wire n672;
   wire n739;
   wire n902;
   wire n925;
   wire n984;
   wire n989;
   wire n1060;
   wire n1061;
   wire n1102;
   wire n1251;
   wire n1495;
   wire n1501;
   wire n1502;
   wire n1503;
   wire n1504;
   wire n1505;
   wire n1506;
   wire n1507;
   wire n1508;
   wire n1509;
   wire n1510;
   wire n1511;
   wire n1512;
   wire n1513;
   wire n1514;
   wire n1515;
   wire n1516;
   wire n1517;
   wire n1518;
   wire n1519;
   wire n1520;
   wire n1521;
   wire n1522;
   wire n1523;
   wire n1524;
   wire n1525;
   wire n1526;
   wire n1527;
   wire n1528;
   wire n1529;
   wire n1530;
   wire n1531;
   wire n1532;
   wire n1533;
   wire n1534;
   wire n1535;
   wire n1536;
   wire n1537;
   wire n1538;
   wire n1539;
   wire n1540;
   wire n1541;
   wire n1542;
   wire n1543;
   wire n1544;
   wire n1545;
   wire n1546;
   wire n1547;
   wire n1548;
   wire n1549;
   wire n1550;
   wire n1551;
   wire n1552;
   wire n1553;
   wire n1554;
   wire n1555;
   wire n1556;
   wire n1557;
   wire n1558;
   wire n1559;
   wire n1560;
   wire n1561;
   wire n1562;
   wire n1563;
   wire n1564;
   wire n1565;
   wire n1566;
   wire n1567;
   wire n1568;
   wire n1569;
   wire n1570;
   wire n1571;
   wire n1572;
   wire n1573;
   wire n1574;
   wire n1575;
   wire n1576;
   wire n1577;
   wire n1578;
   wire n1579;
   wire n1580;
   wire n1581;
   wire n1582;
   wire n1583;
   wire n1584;
   wire n1585;
   wire n1586;
   wire n1587;
   wire n1588;
   wire n1589;
   wire n1590;
   wire n1591;
   wire n1592;
   wire n1593;
   wire n1594;
   wire n1595;
   wire n1596;
   wire n1597;
   wire n1598;
   wire n1599;
   wire n1600;

   OAI32X1 U1 (.Y(n766), 
	.B1(n767), 
	.B0(n121), 
	.A2(n576), 
	.A1(sboxw[26]), 
	.A0(n730));
   AOI31X1 U2 (.Y(n735), 
	.B0(n742), 
	.A2(n1578), 
	.A1(n616), 
	.A0(sboxw[28]));
   OAI31X1 U3 (.Y(n640), 
	.B0(n641), 
	.A2(sboxw[26]), 
	.A1(sboxw[28]), 
	.A0(n616));
   OAI222XL U4 (.Y(n1318), 
	.C1(n230), 
	.C0(n1321), 
	.B1(n24), 
	.B0(n246), 
	.A1(n25), 
	.A0(n243));
   AOI222X1 U5 (.Y(n1300), 
	.C1(n55), 
	.C0(n1503), 
	.B1(n239), 
	.B0(n24), 
	.A1(n635), 
	.A0(n247));
   NAND2X1 U6 (.Y(n240), 
	.B(n23), 
	.A(n247));
   NAND2X1 U7 (.Y(n1), 
	.B(n204), 
	.A(sboxw[18]));
   NAND2X1 U8 (.Y(n2), 
	.B(n1592), 
	.A(sboxw[28]));
   NAND2X1 U9 (.Y(n3), 
	.B(n1552), 
	.A(sboxw[2]));
   NAND2X1 U10 (.Y(n4), 
	.B(n1594), 
	.A(n1592));
   NAND2X1 U11 (.Y(n5), 
	.B(n170), 
	.A(n167));
   NAND2X1 U12 (.Y(n6), 
	.B(n151), 
	.A(n148));
   NAND2X1 U13 (.Y(n7), 
	.B(n170), 
	.A(n166));
   NAND2X1 U14 (.Y(n8), 
	.B(n151), 
	.A(n147));
   NAND2X1 U15 (.Y(n9), 
	.B(n1545), 
	.A(sboxw[3]));
   NAND2X1 U16 (.Y(n10), 
	.B(n139), 
	.A(n136));
   NAND2X1 U17 (.Y(n11), 
	.B(n139), 
	.A(n135));
   NAND2X1 U18 (.Y(n12), 
	.B(sboxw[10]), 
	.A(n60));
   NAND2X1 U19 (.Y(n13), 
	.B(n1251), 
	.A(n1511));
   NAND2X1 U20 (.Y(n14), 
	.B(n63), 
	.A(sboxw[26]));
   NAND2X1 U21 (.Y(n15), 
	.B(n197), 
	.A(n207));
   NAND2X1 U22 (.Y(n16), 
	.B(n1545), 
	.A(n1555));
   NAND2X1 U23 (.Y(n17), 
	.B(sboxw[10]), 
	.A(n1507));
   NAND2X1 U24 (.Y(n18), 
	.B(n56), 
	.A(sboxw[18]));
   NAND2X1 U25 (.Y(n19), 
	.B(n57), 
	.A(sboxw[2]));
   NAND2X1 U26 (.Y(n20), 
	.B(n207), 
	.A(sboxw[20]));
   NAND2X1 U27 (.Y(n21), 
	.B(n1555), 
	.A(sboxw[4]));
   NAND2X1 U28 (.Y(n22), 
	.B(sboxw[27]), 
	.A(sboxw[28]));
   INVX1 U29 (.Y(n247), 
	.A(n55));
   OAI31X1 U30 (.Y(n411), 
	.B0(n412), 
	.A2(sboxw[2]), 
	.A1(sboxw[4]), 
	.A0(n387));
   INVX1 U31 (.Y(n616), 
	.A(n32));
   OAI31X1 U32 (.Y(n994), 
	.B0(n995), 
	.A2(sboxw[18]), 
	.A1(sboxw[20]), 
	.A0(n970));
   INVX1 U33 (.Y(n970), 
	.A(n33));
   INVX1 U34 (.Y(n387), 
	.A(n34));
   INVX1 U35 (.Y(n23), 
	.A(n54));
   OAI222XL U36 (.Y(n1392), 
	.C1(n25), 
	.C0(n242), 
	.B1(n1394), 
	.B0(n23), 
	.A1(n1517), 
	.A0(n1374));
   INVX1 U37 (.Y(n576), 
	.A(n26));
   AOI22XL U38 (.Y(n587), 
	.B1(n616), 
	.B0(n1583), 
	.A1(sboxw[26]), 
	.A0(n123));
   INVX1 U39 (.Y(n24), 
	.A(n65));
   OAI32X1 U40 (.Y(n504), 
	.B1(n505), 
	.B0(n7), 
	.A2(n347), 
	.A1(sboxw[2]), 
	.A0(n468));
   INVX1 U41 (.Y(n347), 
	.A(n28));
   OAI32X1 U42 (.Y(n1087), 
	.B1(n1088), 
	.B0(n118), 
	.A2(n930), 
	.A1(sboxw[18]), 
	.A0(n1051));
   INVX1 U43 (.Y(n930), 
	.A(n27));
   AOI22XL U44 (.Y(n358), 
	.B1(n387), 
	.B0(n1559), 
	.A1(sboxw[2]), 
	.A0(n117));
   AOI22XL U45 (.Y(n941), 
	.B1(n970), 
	.B0(n211), 
	.A1(sboxw[18]), 
	.A0(n120));
   INVX1 U46 (.Y(n25), 
	.A(n50));
   AOI222X1 U57 (.Y(n799), 
	.C1(n26), 
	.C0(n1575), 
	.B1(n122), 
	.B0(n1574), 
	.A1(n121), 
	.A0(n1582));
   AOI222X1 U58 (.Y(n1148), 
	.C1(n27), 
	.C0(n190), 
	.B1(n119), 
	.B0(n198), 
	.A1(n8), 
	.A0(n187));
   AOI222X1 U59 (.Y(n537), 
	.C1(n28), 
	.C0(n1538), 
	.B1(n116), 
	.B0(n1546), 
	.A1(n115), 
	.A0(n1534));
   NAND2X1 U60 (.Y(n1069), 
	.B(n29), 
	.A(n202));
   NAND2X1 U61 (.Y(n486), 
	.B(n31), 
	.A(n1550));
   INVX1 U62 (.Y(n1579), 
	.A(n602));
   INVX1 U63 (.Y(n179), 
	.A(n956));
   INVX1 U64 (.Y(n1526), 
	.A(n373));
   AOI21X1 U65 (.Y(n825), 
	.B0(n668), 
	.A1(n1574), 
	.A0(n121));
   AOI21X1 U66 (.Y(n1174), 
	.B0(n1022), 
	.A1(n198), 
	.A0(n118));
   AOI21X1 U67 (.Y(n682), 
	.B0(n439), 
	.A1(n1546), 
	.A0(n115));
   NAND2X1 U68 (.Y(n964), 
	.B(n29), 
	.A(n180));
   NAND2X1 U69 (.Y(n381), 
	.B(n31), 
	.A(n1527));
   AND2X2 U70 (.Y(n26), 
	.B(n10), 
	.A(n123));
   AND2X2 U71 (.Y(n27), 
	.B(n6), 
	.A(n120));
   AND2X2 U72 (.Y(n28), 
	.B(n5), 
	.A(n117));
   INVX1 U73 (.Y(n125), 
	.A(n126));
   INVX1 U74 (.Y(n123), 
	.A(n30));
   INVX1 U75 (.Y(n120), 
	.A(n29));
   INVX1 U76 (.Y(n117), 
	.A(n31));
   INVX1 U80 (.Y(n127), 
	.A(n125));
   NAND2X1 U81 (.Y(n748), 
	.B(n30), 
	.A(n1576));
   INVX1 U82 (.Y(n273), 
	.A(n1265));
   NAND2X1 U83 (.Y(n610), 
	.B(n30), 
	.A(n1580));
   AND2X2 U84 (.Y(n29), 
	.B(n147), 
	.A(n150));
   AND2X2 U85 (.Y(n30), 
	.B(n135), 
	.A(sboxw[24]));
   AND2X2 U86 (.Y(n31), 
	.B(n166), 
	.A(sboxw[0]));
   OAI21XL U87 (.Y(n1053), 
	.B0(n1054), 
	.A1(n985), 
	.A0(n36));
   OAI21XL U88 (.Y(n470), 
	.B0(n471), 
	.A1(n402), 
	.A0(n37));
   INVX1 U89 (.Y(n1565), 
	.A(n652));
   INVX1 U90 (.Y(n194), 
	.A(n1006));
   INVX1 U91 (.Y(n1542), 
	.A(n423));
   INVX1 U93 (.Y(n190), 
	.A(n937));
   INVX1 U94 (.Y(n635), 
	.A(n1374));
   INVX1 U95 (.Y(n1495), 
	.A(n1311));
   NOR2X1 U96 (.Y(n668), 
	.B(n11), 
	.A(n814));
   NOR2X1 U97 (.Y(n1022), 
	.B(n8), 
	.A(n1163));
   NOR2X1 U98 (.Y(n439), 
	.B(n7), 
	.A(n552));
   OAI221XL U99 (.Y(n1193), 
	.C0(n955), 
	.B1(n1194), 
	.B0(n930), 
	.A1(n954), 
	.A0(n27));
   OAI221XL U100 (.Y(n701), 
	.C0(n372), 
	.B1(n702), 
	.B0(n347), 
	.A1(n371), 
	.A0(n28));
   NOR2X1 U101 (.Y(n313), 
	.B(n125), 
	.A(n1290));
   NAND2X1 U102 (.Y(n1384), 
	.B(n1495), 
	.A(n65));
   NOR2X1 U103 (.Y(n627), 
	.B(n26), 
	.A(n583));
   NOR2X1 U104 (.Y(n981), 
	.B(n27), 
	.A(n937));
   NOR2X1 U105 (.Y(n398), 
	.B(n28), 
	.A(n354));
   NOR2X1 U106 (.Y(n1287), 
	.B(n153), 
	.A(n54));
   NOR2X1 U107 (.Y(n933), 
	.B(n143), 
	.A(n36));
   NOR2X1 U108 (.Y(n350), 
	.B(sboxw[5]), 
	.A(n37));
   AOI31X1 U109 (.Y(n592), 
	.B0(n599), 
	.A2(n575), 
	.A1(n598), 
	.A0(n597));
   AOI31X1 U110 (.Y(n946), 
	.B0(n953), 
	.A2(n929), 
	.A1(n952), 
	.A0(n951));
   AOI31X1 U111 (.Y(n363), 
	.B0(n370), 
	.A2(n346), 
	.A1(n369), 
	.A0(n368));
   AOI31X1 U112 (.Y(n593), 
	.B0(n130), 
	.A2(n596), 
	.A1(n595), 
	.A0(n594));
   AOI31X1 U113 (.Y(n947), 
	.B0(sboxw[21]), 
	.A2(n950), 
	.A1(n949), 
	.A0(n948));
   AOI31X1 U114 (.Y(n364), 
	.B0(n159), 
	.A2(n367), 
	.A1(n366), 
	.A0(n365));
   NOR2X1 U115 (.Y(n921), 
	.B(n146), 
	.A(n1163));
   NOR2X1 U116 (.Y(n338), 
	.B(n167), 
	.A(n552));
   INVX1 U117 (.Y(n1578), 
	.A(n604));
   INVX1 U118 (.Y(n185), 
	.A(n958));
   INVX1 U119 (.Y(n1532), 
	.A(n375));
   INVX1 U120 (.Y(n413), 
	.A(n1342));
   NAND2X1 U121 (.Y(n959), 
	.B(n196), 
	.A(n38));
   NAND2X1 U122 (.Y(n376), 
	.B(n1544), 
	.A(n39));
   INVX1 U123 (.Y(n1577), 
	.A(n845));
   INVX1 U124 (.Y(n1531), 
	.A(n702));
   INVX1 U125 (.Y(n184), 
	.A(n1194));
   NAND2X1 U126 (.Y(n602), 
	.B(n1581), 
	.A(n1591));
   NAND2X1 U127 (.Y(n956), 
	.B(n181), 
	.A(n196));
   NAND2X1 U128 (.Y(n373), 
	.B(n1528), 
	.A(n1544));
   INVX1 U129 (.Y(n150), 
	.A(n151));
   INVX1 U130 (.Y(n135), 
	.A(n136));
   INVX1 U131 (.Y(n147), 
	.A(n146));
   INVX1 U132 (.Y(n166), 
	.A(n167));
   OAI21XL U133 (.Y(n732), 
	.B0(n733), 
	.A1(n631), 
	.A0(n35));
   INVX1 U134 (.Y(n1060), 
	.A(n1327));
   INVX1 U135 (.Y(n406), 
	.A(n323));
   INVX1 U136 (.Y(n1580), 
	.A(n881));
   INVX1 U137 (.Y(n180), 
	.A(n1230));
   INVX1 U138 (.Y(n1527), 
	.A(n1474));
   INVX1 U139 (.Y(n925), 
	.A(n1371));
   INVX1 U140 (.Y(n153), 
	.A(sboxw[13]));
   AND2X2 U141 (.Y(n32), 
	.B(n136), 
	.A(sboxw[24]));
   AND2X2 U142 (.Y(n33), 
	.B(n146), 
	.A(n150));
   AND2X2 U143 (.Y(n34), 
	.B(n167), 
	.A(sboxw[0]));
   INVX1 U144 (.Y(n129), 
	.A(n131));
   INVX1 U145 (.Y(n142), 
	.A(sboxw[21]));
   INVX1 U146 (.Y(n161), 
	.A(n162));
   INVX1 U148 (.Y(n1503), 
	.A(n1308));
   INVX1 U149 (.Y(n1581), 
	.A(n599));
   INVX1 U150 (.Y(n181), 
	.A(n953));
   INVX1 U151 (.Y(n1528), 
	.A(n370));
   INVX1 U152 (.Y(n1582), 
	.A(n814));
   INVX1 U153 (.Y(n739), 
	.A(n1290));
   INVX1 U155 (.Y(n1575), 
	.A(n583));
   INVX1 U157 (.Y(n1538), 
	.A(n354));
   INVX1 U158 (.Y(n187), 
	.A(n1163));
   INVX1 U159 (.Y(n1534), 
	.A(n552));
   AND2X2 U160 (.Y(n35), 
	.B(n139), 
	.A(n135));
   INVX1 U161 (.Y(n121), 
	.A(n35));
   AND2X2 U162 (.Y(n36), 
	.B(n151), 
	.A(n147));
   INVX1 U163 (.Y(n118), 
	.A(n36));
   AND2X2 U164 (.Y(n37), 
	.B(n170), 
	.A(n166));
   INVX1 U165 (.Y(n115), 
	.A(n37));
   INVX1 U166 (.Y(n126), 
	.A(n240));
   OAI221XL U167 (.Y(n844), 
	.C0(n601), 
	.B1(n845), 
	.B0(n576), 
	.A1(n600), 
	.A0(n26));
   NOR2X1 U168 (.Y(n579), 
	.B(n130), 
	.A(n35));
   NOR2X1 U169 (.Y(n567), 
	.B(n136), 
	.A(n814));
   NAND2X1 U170 (.Y(n605), 
	.B(n1591), 
	.A(n40));
   NAND2X1 U171 (.Y(n1265), 
	.B(n1102), 
	.A(n49));
   OAI21XL U172 (.Y(n591), 
	.B0(n601), 
	.A1(n600), 
	.A0(n135));
   OAI21XL U173 (.Y(n945), 
	.B0(n955), 
	.A1(n954), 
	.A0(n147));
   OAI21XL U174 (.Y(n362), 
	.B0(n372), 
	.A1(n371), 
	.A0(n166));
   NAND2X1 U175 (.Y(n1296), 
	.B(n65), 
	.A(n276));
   INVX1 U176 (.Y(n276), 
	.A(n282));
   INVX1 U178 (.Y(n1574), 
	.A(n631));
   INVX1 U180 (.Y(n1546), 
	.A(n402));
   INVX1 U182 (.Y(n198), 
	.A(n985));
   INVX1 U183 (.Y(n1560), 
	.A(n597));
   INVX1 U184 (.Y(n186), 
	.A(n951));
   INVX1 U185 (.Y(n1533), 
	.A(n368));
   INVX1 U186 (.Y(n1576), 
	.A(n767));
   INVX1 U187 (.Y(n202), 
	.A(n1088));
   INVX1 U188 (.Y(n1550), 
	.A(n505));
   INVX1 U191 (.Y(n229), 
	.A(n1414));
   AND2X2 U192 (.Y(n38), 
	.B(n151), 
	.A(n148));
   INVX1 U193 (.Y(n119), 
	.A(n38));
   AND2X2 U194 (.Y(n39), 
	.B(n170), 
	.A(n167));
   INVX1 U195 (.Y(n116), 
	.A(n39));
   AND2X2 U196 (.Y(n40), 
	.B(n139), 
	.A(n136));
   INVX1 U197 (.Y(n122), 
	.A(n40));
   INVX1 U203 (.Y(n1591), 
	.A(n4));
   INVX1 U204 (.Y(n196), 
	.A(n15));
   INVX1 U205 (.Y(n1544), 
	.A(n16));
   OAI222XL U206 (.Y(n1083), 
	.C1(n1096), 
	.C0(n143), 
	.B1(n958), 
	.B0(n1095), 
	.A1(n142), 
	.A0(n1094));
   AOI21X1 U207 (.Y(n1095), 
	.B0(n186), 
	.A1(n6), 
	.A0(n196));
   AOI221X1 U208 (.Y(n1094), 
	.C0(n1100), 
	.B1(n56), 
	.B0(n33), 
	.A1(n38), 
	.A0(n205));
   AOI211X1 U209 (.Y(n1096), 
	.C0(n1098), 
	.B0(n1097), 
	.A1(n146), 
	.A0(n190));
   OAI222XL U210 (.Y(n500), 
	.C1(n513), 
	.C0(n159), 
	.B1(n375), 
	.B0(n512), 
	.A1(n163), 
	.A0(n511));
   AOI21X1 U211 (.Y(n512), 
	.B0(n1533), 
	.A1(n5), 
	.A0(n1544));
   AOI221X1 U212 (.Y(n511), 
	.C0(n517), 
	.B1(n57), 
	.B0(n34), 
	.A1(n39), 
	.A0(n1553));
   AOI211X1 U213 (.Y(n513), 
	.C0(n515), 
	.B0(n514), 
	.A1(n167), 
	.A0(n1538));
   OAI211X1 U214 (.Y(n880), 
	.C0(n883), 
	.B0(n882), 
	.A1(n881), 
	.A0(n26));
   AOI31X1 U215 (.Y(n882), 
	.B0(n1570), 
	.A2(n577), 
	.A1(n730), 
	.A0(n26));
   AOI222X1 U216 (.Y(n883), 
	.C1(n616), 
	.C0(n1579), 
	.B1(n122), 
	.B0(n1573), 
	.A1(n884), 
	.A0(sboxw[29]));
   INVX1 U217 (.Y(n1570), 
	.A(n837));
   OAI211X1 U218 (.Y(n1473), 
	.C0(n1476), 
	.B0(n1475), 
	.A1(n1474), 
	.A0(n28));
   AOI31X1 U219 (.Y(n1475), 
	.B0(n1530), 
	.A2(n348), 
	.A1(n468), 
	.A0(n28));
   AOI222X1 U220 (.Y(n1476), 
	.C1(n387), 
	.C0(n1526), 
	.B1(n5), 
	.B0(n1525), 
	.A1(n1477), 
	.A0(sboxw[5]));
   INVX1 U221 (.Y(n1530), 
	.A(n694));
   OAI221XL U222 (.Y(n1036), 
	.C0(n1050), 
	.B1(n142), 
	.B0(n1049), 
	.A1(n953), 
	.A0(n1048));
   AOI222X1 U223 (.Y(n1048), 
	.C1(n196), 
	.C0(n36), 
	.B1(n204), 
	.B0(n29), 
	.A1(n970), 
	.A0(n56));
   AOI32X1 U224 (.Y(n1050), 
	.B1(sboxw[16]), 
	.B0(n178), 
	.A2(n931), 
	.A1(n120), 
	.A0(n1051));
   AOI211X1 U225 (.Y(n1049), 
	.C0(n1053), 
	.B0(n1052), 
	.A1(n147), 
	.A0(n190));
   OAI221XL U226 (.Y(n453), 
	.C0(n467), 
	.B1(n163), 
	.B0(n466), 
	.A1(n370), 
	.A0(n465));
   AOI222X1 U227 (.Y(n465), 
	.C1(n1544), 
	.C0(n37), 
	.B1(n1552), 
	.B0(n31), 
	.A1(n387), 
	.A0(n57));
   AOI32X1 U228 (.Y(n467), 
	.B1(sboxw[0]), 
	.B0(n1525), 
	.A2(n348), 
	.A1(n117), 
	.A0(n468));
   AOI211X1 U229 (.Y(n466), 
	.C0(n470), 
	.B0(n469), 
	.A1(sboxw[1]), 
	.A0(n1538));
   AOI211X1 U230 (.Y(n800), 
	.C0(n1569), 
	.B0(n606), 
	.A1(n616), 
	.A0(n566));
   INVX1 U231 (.Y(n1569), 
	.A(n717));
   AOI211X1 U232 (.Y(n1149), 
	.C0(n192), 
	.B0(n960), 
	.A1(n970), 
	.A0(n920));
   INVX1 U233 (.Y(n192), 
	.A(n1038));
   AOI211X1 U234 (.Y(n538), 
	.C0(n1540), 
	.B0(n377), 
	.A1(n387), 
	.A0(n337));
   INVX1 U235 (.Y(n1540), 
	.A(n455));
   NAND2X1 U236 (.Y(n937), 
	.B(n211), 
	.A(n196));
   OAI211X1 U237 (.Y(n1229), 
	.C0(n1232), 
	.B0(n1231), 
	.A1(n1230), 
	.A0(n27));
   AOI31X1 U238 (.Y(n1231), 
	.B0(n183), 
	.A2(n931), 
	.A1(n1051), 
	.A0(n27));
   AOI222X1 U239 (.Y(n1232), 
	.C1(n970), 
	.C0(n179), 
	.B1(n6), 
	.B0(n178), 
	.A1(n1233), 
	.A0(sboxw[21]));
   INVX1 U240 (.Y(n183), 
	.A(n1186));
   NOR2X1 U241 (.Y(n1178), 
	.B(n190), 
	.A(n199));
   AOI211X1 U242 (.Y(n1074), 
	.C0(n193), 
	.B0(n960), 
	.A1(n119), 
	.A0(n203));
   INVX1 U243 (.Y(n193), 
	.A(n1081));
   AOI22X1 U244 (.Y(n826), 
	.B1(n1586), 
	.B0(n11), 
	.A1(n1585), 
	.A0(n135));
   AOI22X1 U245 (.Y(n1175), 
	.B1(n61), 
	.B0(n118), 
	.A1(n195), 
	.A0(n147));
   AOI22X1 U246 (.Y(n683), 
	.B1(n62), 
	.B0(n115), 
	.A1(n1543), 
	.A0(n166));
   NAND2X1 U247 (.Y(n1081), 
	.B(n151), 
	.A(n195));
   NAND2X1 U248 (.Y(n498), 
	.B(n169), 
	.A(n1543));
   NAND2X1 U249 (.Y(n717), 
	.B(n123), 
	.A(n1585));
   NAND2X1 U250 (.Y(n1038), 
	.B(n120), 
	.A(n195));
   NAND2X1 U251 (.Y(n455), 
	.B(n117), 
	.A(n1543));
   NAND2X1 U252 (.Y(n733), 
	.B(n1585), 
	.A(n35));
   NAND2X1 U253 (.Y(n1054), 
	.B(n195), 
	.A(n36));
   NAND2X1 U254 (.Y(n471), 
	.B(n1543), 
	.A(n37));
   AOI21X1 U255 (.Y(n968), 
	.B0(n1190), 
	.A1(n195), 
	.A0(n119));
   NAND4BXL U256 (.Y(n784), 
	.D(n797), 
	.C(n796), 
	.B(n610), 
	.AN(n795));
   AOI22X1 U257 (.Y(n796), 
	.B1(n63), 
	.B0(n579), 
	.A1(n32), 
	.A0(n801));
   AOI211X1 U258 (.Y(n797), 
	.C0(n725), 
	.B0(n798), 
	.A1(sboxw[25]), 
	.A0(n789));
   AOI21X1 U259 (.Y(n798), 
	.B0(n129), 
	.A1(n800), 
	.A0(n799));
   NAND4BXL U260 (.Y(n1133), 
	.D(n1146), 
	.C(n1145), 
	.B(n964), 
	.AN(n1144));
   AOI22X1 U261 (.Y(n1145), 
	.B1(n64), 
	.B0(n933), 
	.A1(n33), 
	.A0(n1150));
   AOI211X1 U262 (.Y(n1146), 
	.C0(n1046), 
	.B0(n1147), 
	.A1(sboxw[17]), 
	.A0(n1138));
   AOI21X1 U263 (.Y(n1147), 
	.B0(n142), 
	.A1(n1149), 
	.A0(n1148));
   NAND4BXL U264 (.Y(n522), 
	.D(n535), 
	.C(n534), 
	.B(n381), 
	.AN(n533));
   AOI22X1 U265 (.Y(n534), 
	.B1(n1536), 
	.B0(n350), 
	.A1(n34), 
	.A0(n539));
   AOI211X1 U266 (.Y(n535), 
	.C0(n463), 
	.B0(n536), 
	.A1(sboxw[1]), 
	.A0(n527));
   AOI21X1 U267 (.Y(n536), 
	.B0(n161), 
	.A1(n538), 
	.A0(n537));
   NAND4BXL U268 (.Y(n1097), 
	.D(n1090), 
	.C(n1081), 
	.B(n927), 
	.AN(n1099));
   NAND4BXL U269 (.Y(n514), 
	.D(n507), 
	.C(n498), 
	.B(n344), 
	.AN(n516));
   NAND4X1 U270 (.Y(n884), 
	.D(n886), 
	.C(n885), 
	.B(n769), 
	.A(n846));
   AOI222X1 U271 (.Y(n886), 
	.C1(n616), 
	.C0(n1586), 
	.B1(n123), 
	.B0(n1575), 
	.A1(n121), 
	.A0(n67));
   AOI21X1 U272 (.Y(n885), 
	.B0(n1565), 
	.A1(n40), 
	.A0(n1574));
   NAND4X1 U273 (.Y(n1233), 
	.D(n1235), 
	.C(n1234), 
	.B(n1090), 
	.A(n1195));
   AOI222X1 U274 (.Y(n1235), 
	.C1(n970), 
	.C0(n61), 
	.B1(n120), 
	.B0(n190), 
	.A1(n8), 
	.A0(n199));
   AOI21X1 U275 (.Y(n1234), 
	.B0(n194), 
	.A1(n38), 
	.A0(n198));
   NAND4X1 U276 (.Y(n1477), 
	.D(n1479), 
	.C(n1478), 
	.B(n507), 
	.A(n703));
   AOI222X1 U277 (.Y(n1479), 
	.C1(n387), 
	.C0(n62), 
	.B1(n117), 
	.B0(n1538), 
	.A1(n7), 
	.A0(n1547));
   AOI21X1 U278 (.Y(n1478), 
	.B0(n1542), 
	.A1(n39), 
	.A0(n1546));
   NAND2X1 U279 (.Y(n652), 
	.B(n26), 
	.A(n1585));
   NAND2X1 U280 (.Y(n1006), 
	.B(n27), 
	.A(n195));
   NAND2X1 U281 (.Y(n423), 
	.B(n28), 
	.A(n1543));
   OAI21XL U282 (.Y(n1177), 
	.B0(n1179), 
	.A1(n970), 
	.A0(n1178));
   AOI31X1 U283 (.Y(n926), 
	.B0(n142), 
	.A2(n928), 
	.A1(n200), 
	.A0(n927));
   AOI21X1 U284 (.Y(n928), 
	.B0(n201), 
	.A1(n147), 
	.A0(n195));
   INVX1 U285 (.Y(n201), 
	.A(n929));
   AOI31X1 U286 (.Y(n343), 
	.B0(n161), 
	.A2(n345), 
	.A1(n1548), 
	.A0(n344));
   AOI21X1 U287 (.Y(n345), 
	.B0(n1549), 
	.A1(n166), 
	.A0(n1543));
   INVX1 U288 (.Y(n1549), 
	.A(n346));
   NOR2X1 U289 (.Y(n291), 
	.B(n153), 
	.A(n1515));
   NAND2X1 U290 (.Y(n1308), 
	.B(n1515), 
	.A(n1507));
   NAND2X1 U291 (.Y(n814), 
	.B(n1583), 
	.A(n63));
   NAND2X1 U292 (.Y(n1163), 
	.B(n211), 
	.A(n64));
   NAND2X1 U293 (.Y(n552), 
	.B(n1559), 
	.A(n1536));
   AOI222X1 U294 (.Y(n261), 
	.C1(n1502), 
	.C0(n65), 
	.B1(n1495), 
	.B0(n50), 
	.A1(n125), 
	.A0(n58));
   NAND2X1 U295 (.Y(n599), 
	.B(n129), 
	.A(n1583));
   NAND2X1 U296 (.Y(n953), 
	.B(n142), 
	.A(n211));
   NAND2X1 U297 (.Y(n370), 
	.B(n161), 
	.A(n1559));
   NAND2X1 U298 (.Y(n1342), 
	.B(n1515), 
	.A(n153));
   NAND2X1 U299 (.Y(n1290), 
	.B(n1515), 
	.A(n1102));
   NAND2X1 U300 (.Y(n604), 
	.B(n1583), 
	.A(n130));
   NAND2X1 U301 (.Y(n958), 
	.B(n211), 
	.A(sboxw[21]));
   NAND2X1 U302 (.Y(n375), 
	.B(n1559), 
	.A(n162));
   OAI222XL U303 (.Y(n590), 
	.C1(n605), 
	.C0(n604), 
	.B1(n128), 
	.B0(n603), 
	.A1(n602), 
	.A0(n26));
   AOI211X1 U304 (.Y(n603), 
	.C0(n589), 
	.B0(n606), 
	.A1(n123), 
	.A0(n63));
   OAI222XL U305 (.Y(n944), 
	.C1(n959), 
	.C0(n958), 
	.B1(n142), 
	.B0(n957), 
	.A1(n956), 
	.A0(n27));
   AOI211X1 U306 (.Y(n957), 
	.C0(n943), 
	.B0(n960), 
	.A1(n120), 
	.A0(n64));
   OAI222XL U307 (.Y(n361), 
	.C1(n376), 
	.C0(n375), 
	.B1(n163), 
	.B0(n374), 
	.A1(n373), 
	.A0(n28));
   AOI211X1 U308 (.Y(n374), 
	.C0(n360), 
	.B0(n377), 
	.A1(n117), 
	.A0(n1536));
   AOI222XL U309 (.Y(n1418), 
	.C1(n25), 
	.C0(n1503), 
	.B1(n125), 
	.B0(n739), 
	.A1(n54), 
	.A0(n1506));
   OAI32X1 U310 (.Y(n1255), 
	.B1(n954), 
	.B0(n33), 
	.A2(n142), 
	.A1(n1256), 
	.A0(n211));
   AOI21X1 U311 (.Y(n1256), 
	.B0(n38), 
	.A1(n118), 
	.A0(n1051));
   OAI32X1 U312 (.Y(n1499), 
	.B1(n371), 
	.B0(n34), 
	.A2(n163), 
	.A1(n1500), 
	.A0(n1559));
   AOI21X1 U313 (.Y(n1500), 
	.B0(n39), 
	.A1(n7), 
	.A0(n468));
   NAND2X1 U314 (.Y(n1311), 
	.B(n1515), 
	.A(n60));
   OAI222XL U315 (.Y(n762), 
	.C1(n775), 
	.C0(sboxw[29]), 
	.B1(n604), 
	.B0(n774), 
	.A1(n128), 
	.A0(n773));
   AOI21X1 U316 (.Y(n774), 
	.B0(n1560), 
	.A1(n10), 
	.A0(n1591));
   AOI221X1 U317 (.Y(n773), 
	.C0(n779), 
	.B1(n1593), 
	.B0(n32), 
	.A1(n40), 
	.A0(n1588));
   AOI211X1 U318 (.Y(n775), 
	.C0(n777), 
	.B0(n776), 
	.A1(n136), 
	.A0(n1575));
   NAND2X1 U319 (.Y(n1374), 
	.B(n1515), 
	.A(n58));
   NAND2X1 U320 (.Y(n769), 
	.B(n66), 
	.A(n35));
   NAND2X1 U321 (.Y(n1090), 
	.B(n203), 
	.A(n36));
   NAND2X1 U322 (.Y(n507), 
	.B(n1551), 
	.A(n37));
   NAND2X1 U323 (.Y(n249), 
	.B(n124), 
	.A(n1502));
   NAND2X1 U324 (.Y(n1284), 
	.B(n1517), 
	.A(n1506));
   NOR3X1 U325 (.Y(n1286), 
	.C(n1342), 
	.B(n65), 
	.A(n13));
   NOR3X1 U326 (.Y(n932), 
	.C(n15), 
	.B(n29), 
	.A(n958));
   NOR3X1 U327 (.Y(n349), 
	.C(n16), 
	.B(n31), 
	.A(n375));
   NAND2X1 U328 (.Y(n583), 
	.B(n1583), 
	.A(n1591));
   NAND2X1 U329 (.Y(n354), 
	.B(n1559), 
	.A(n1544));
   NOR2X1 U330 (.Y(n829), 
	.B(n1575), 
	.A(n67));
   NOR2X1 U331 (.Y(n686), 
	.B(n1538), 
	.A(n1547));
   NAND2X1 U332 (.Y(n718), 
	.B(n26), 
	.A(n67));
   NAND2X1 U333 (.Y(n1039), 
	.B(n27), 
	.A(n199));
   NAND2X1 U334 (.Y(n456), 
	.B(n28), 
	.A(n1547));
   OAI221XL U335 (.Y(n715), 
	.C0(n729), 
	.B1(n128), 
	.B0(n728), 
	.A1(n599), 
	.A0(n727));
   AOI32X1 U336 (.Y(n729), 
	.B1(sboxw[24]), 
	.B0(n1573), 
	.A2(n577), 
	.A1(n123), 
	.A0(n730));
   AOI222X1 U337 (.Y(n727), 
	.C1(n1591), 
	.C0(n35), 
	.B1(n1590), 
	.B0(n30), 
	.A1(n616), 
	.A0(n1593));
   AOI211X1 U338 (.Y(n728), 
	.C0(n732), 
	.B0(n731), 
	.A1(n135), 
	.A0(n1575));
   AOI211X1 U339 (.Y(n753), 
	.C0(n1584), 
	.B0(n606), 
	.A1(n10), 
	.A0(n66));
   INVX1 U340 (.Y(n1584), 
	.A(n760));
   AOI211X1 U341 (.Y(n491), 
	.C0(n1541), 
	.B0(n377), 
	.A1(n116), 
	.A0(n1551));
   INVX1 U342 (.Y(n1541), 
	.A(n498));
   NAND2X1 U343 (.Y(n248), 
	.B(n125), 
	.A(n1506));
   INVX1 U344 (.Y(n200), 
	.A(n1190));
   INVX1 U345 (.Y(n1548), 
	.A(n698));
   NAND2X1 U346 (.Y(n598), 
	.B(n1593), 
	.A(n26));
   NAND2X1 U347 (.Y(n952), 
	.B(n56), 
	.A(n27));
   NAND2X1 U348 (.Y(n369), 
	.B(n57), 
	.A(n28));
   OAI211X1 U349 (.Y(n646), 
	.C0(n595), 
	.B0(n647), 
	.A1(n135), 
	.A0(n4));
   OAI211X1 U350 (.Y(n1000), 
	.C0(n949), 
	.B0(n1001), 
	.A1(sboxw[17]), 
	.A0(n15));
   OAI211X1 U351 (.Y(n417), 
	.C0(n366), 
	.B0(n418), 
	.A1(n166), 
	.A0(n16));
   OAI211XL U352 (.Y(n1031), 
	.C0(n927), 
	.B0(n965), 
	.A1(n15), 
	.A0(n930));
   OAI211XL U353 (.Y(n448), 
	.C0(n344), 
	.B0(n382), 
	.A1(n16), 
	.A0(n347));
   OAI211X1 U354 (.Y(n1350), 
	.C0(n1283), 
	.B0(n1298), 
	.A1(n13), 
	.A0(n126));
   NAND2X1 U355 (.Y(n316), 
	.B(n125), 
	.A(n1507));
   NAND2X1 U356 (.Y(n954), 
	.B(n185), 
	.A(n204));
   NAND2X1 U357 (.Y(n371), 
	.B(n1532), 
	.A(n1552));
   NAND2X1 U358 (.Y(n949), 
	.B(n147), 
	.A(n203));
   NAND2X1 U359 (.Y(n366), 
	.B(n166), 
	.A(n1551));
   AOI22X1 U360 (.Y(n615), 
	.B1(n1586), 
	.B0(n576), 
	.A1(n66), 
	.A0(n136));
   AOI22X1 U361 (.Y(n969), 
	.B1(n61), 
	.B0(n930), 
	.A1(n203), 
	.A0(n146));
   AOI22X1 U362 (.Y(n386), 
	.B1(n62), 
	.B0(n347), 
	.A1(n1551), 
	.A0(n167));
   NAND2X1 U363 (.Y(n936), 
	.B(n147), 
	.A(n61));
   NAND2X1 U364 (.Y(n353), 
	.B(n166), 
	.A(n62));
   AOI22X1 U365 (.Y(n647), 
	.B1(n1588), 
	.B0(n32), 
	.A1(n1586), 
	.A0(n121));
   AOI22X1 U366 (.Y(n1001), 
	.B1(n205), 
	.B0(n33), 
	.A1(n61), 
	.A0(n118));
   AOI22X1 U367 (.Y(n418), 
	.B1(n1553), 
	.B0(n34), 
	.A1(n62), 
	.A0(n115));
   AOI31X1 U368 (.Y(n572), 
	.B0(n129), 
	.A2(n574), 
	.A1(n1587), 
	.A0(n573));
   AOI21X1 U369 (.Y(n574), 
	.B0(n1589), 
	.A1(n135), 
	.A0(n1585));
   INVX1 U370 (.Y(n1589), 
	.A(n575));
   NAND2X1 U371 (.Y(n760), 
	.B(n139), 
	.A(n1585));
   NAND2X1 U372 (.Y(n264), 
	.B(n1517), 
	.A(n1061));
   NAND2X1 U373 (.Y(n1055), 
	.B(n150), 
	.A(n64));
   NAND2X1 U374 (.Y(n258), 
	.B(n126), 
	.A(n1506));
   NAND2X1 U375 (.Y(n596), 
	.B(n1585), 
	.A(n32));
   NAND2X1 U376 (.Y(n950), 
	.B(n195), 
	.A(n33));
   NAND2X1 U377 (.Y(n367), 
	.B(n1543), 
	.A(n34));
   NAND2X1 U378 (.Y(n573), 
	.B(n32), 
	.A(n1586));
   NAND2X1 U379 (.Y(n927), 
	.B(n33), 
	.A(n61));
   NAND2X1 U380 (.Y(n344), 
	.B(n34), 
	.A(n62));
   NAND2X1 U381 (.Y(n1283), 
	.B(n59), 
	.A(n55));
   AOI21X1 U382 (.Y(n614), 
	.B0(n841), 
	.A1(n1585), 
	.A0(n122));
   AOI21X1 U383 (.Y(n385), 
	.B0(n698), 
	.A1(n1543), 
	.A0(n116));
   NAND2X1 U384 (.Y(n323), 
	.B(n60), 
	.A(n413));
   OAI22X1 U385 (.Y(n721), 
	.B1(n724), 
	.B0(n130), 
	.A1(n129), 
	.A0(n723));
   AOI21X1 U386 (.Y(n723), 
	.B0(n67), 
	.A1(n138), 
	.A0(n629));
   AOI21X1 U387 (.Y(n724), 
	.B0(n725), 
	.A1(n616), 
	.A0(n63));
   OAI22X1 U388 (.Y(n1042), 
	.B1(n1045), 
	.B0(n143), 
	.A1(n142), 
	.A0(n1044));
   AOI21X1 U389 (.Y(n1044), 
	.B0(n199), 
	.A1(n151), 
	.A0(n983));
   AOI21X1 U390 (.Y(n1045), 
	.B0(n1046), 
	.A1(n970), 
	.A0(n64));
   OAI22X1 U391 (.Y(n459), 
	.B1(n462), 
	.B0(sboxw[5]), 
	.A1(n161), 
	.A0(n461));
   AOI21X1 U392 (.Y(n461), 
	.B0(n1547), 
	.A1(n170), 
	.A0(n400));
   AOI21X1 U393 (.Y(n462), 
	.B0(n463), 
	.A1(n387), 
	.A0(n1536));
   NOR2X1 U394 (.Y(n1240), 
	.B(n33), 
	.A(n46));
   XNOR2X1 U395 (.Y(n46), 
	.B(n150), 
	.A(n211));
   NOR2X1 U396 (.Y(n1484), 
	.B(n34), 
	.A(n47));
   XNOR2X1 U397 (.Y(n47), 
	.B(n168), 
	.A(n1559));
   NAND2X1 U398 (.Y(n881), 
	.B(n1593), 
	.A(n1581));
   NAND2X1 U399 (.Y(n1230), 
	.B(n56), 
	.A(n181));
   NAND2X1 U400 (.Y(n1474), 
	.B(n57), 
	.A(n1528));
   NAND2X1 U401 (.Y(n965), 
	.B(n204), 
	.A(n36));
   NAND2X1 U402 (.Y(n382), 
	.B(n1552), 
	.A(n37));
   NAND2X1 U403 (.Y(n1298), 
	.B(n60), 
	.A(n124));
   AOI22X1 U404 (.Y(n859), 
	.B1(n11), 
	.B0(n1585), 
	.A1(n26), 
	.A0(n1582));
   AOI22X1 U405 (.Y(n1208), 
	.B1(n8), 
	.B0(n195), 
	.A1(n27), 
	.A0(n187));
   AOI22X1 U406 (.Y(n1113), 
	.B1(n7), 
	.B0(n1543), 
	.A1(n28), 
	.A0(n1534));
   NAND2X1 U407 (.Y(n845), 
	.B(n1578), 
	.A(n63));
   NAND2X1 U408 (.Y(n702), 
	.B(n1532), 
	.A(n1536));
   NAND2X1 U409 (.Y(n1194), 
	.B(n185), 
	.A(n64));
   NAND2X1 U410 (.Y(n1186), 
	.B(n147), 
	.A(n1150));
   NAND2X1 U411 (.Y(n694), 
	.B(n166), 
	.A(n539));
   INVX1 U412 (.Y(n1510), 
	.A(n1278));
   NAND2X1 U413 (.Y(n1371), 
	.B(n1061), 
	.A(n54));
   NAND4BXL U414 (.Y(n1407), 
	.D(n249), 
	.C(n264), 
	.B(n1283), 
	.AN(n232));
   NAND4BXL U415 (.Y(n776), 
	.D(n769), 
	.C(n760), 
	.B(n573), 
	.AN(n778));
   NAND4BXL U416 (.Y(n866), 
	.D(n871), 
	.C(n870), 
	.B(n760), 
	.AN(n567));
   AOI222X1 U417 (.Y(n871), 
	.C1(n35), 
	.C0(n1586), 
	.B1(n26), 
	.B0(n1574), 
	.A1(n66), 
	.A0(n40));
   AOI2BB2X1 U418 (.Y(n870), 
	.B1(n137), 
	.B0(n1576), 
	.A1N(n40), 
	.A0N(n829));
   NAND4BXL U419 (.Y(n1215), 
	.D(n1220), 
	.C(n1219), 
	.B(n1081), 
	.AN(n921));
   AOI222X1 U420 (.Y(n1220), 
	.C1(n36), 
	.C0(n61), 
	.B1(n27), 
	.B0(n198), 
	.A1(n203), 
	.A0(n38));
   AOI2BB2X1 U421 (.Y(n1219), 
	.B1(n150), 
	.B0(n202), 
	.A1N(n38), 
	.A0N(n1178));
   NAND4BXL U422 (.Y(n1120), 
	.D(n1125), 
	.C(n1124), 
	.B(n498), 
	.AN(n338));
   AOI222X1 U423 (.Y(n1125), 
	.C1(n37), 
	.C0(n62), 
	.B1(n28), 
	.B0(n1546), 
	.A1(n1551), 
	.A0(n39));
   AOI2BB2X1 U424 (.Y(n1124), 
	.B1(n168), 
	.B0(n1550), 
	.A1N(n39), 
	.A0N(n686));
   NAND2X1 U425 (.Y(n1327), 
	.B(n125), 
	.A(n1061));
   NAND4X1 U426 (.Y(n731), 
	.D(n718), 
	.C(n595), 
	.B(n734), 
	.A(n714));
   NAND4X1 U427 (.Y(n1052), 
	.D(n1039), 
	.C(n949), 
	.B(n1055), 
	.A(n1035));
   NAND4X1 U428 (.Y(n469), 
	.D(n456), 
	.C(n366), 
	.B(n472), 
	.A(n452));
   OAI21XL U429 (.Y(n828), 
	.B0(n830), 
	.A1(n616), 
	.A0(n829));
   OAI21XL U430 (.Y(n685), 
	.B0(n687), 
	.A1(n387), 
	.A0(n686));
   INVX1 U431 (.Y(n178), 
	.A(n1185));
   INVX1 U432 (.Y(n1525), 
	.A(n693));
   NOR2X1 U433 (.Y(n1426), 
	.B(n1061), 
	.A(n1503));
   INVX1 U434 (.Y(n630), 
	.A(n1455));
   AOI221X1 U435 (.Y(n1455), 
	.C0(n303), 
	.B1(n126), 
	.B0(n635), 
	.A1(n55), 
	.A0(n252));
   INVX1 U437 (.Y(n1102), 
	.A(n13));
   AOI221XL U438 (.Y(n1389), 
	.C0(n984), 
	.B1(n25), 
	.B0(n1502), 
	.A1(n124), 
	.A0(n1506));
   INVX1 U439 (.Y(n984), 
	.A(n264));
   INVX1 U440 (.Y(n139), 
	.A(n137));
   INVX1 U441 (.Y(n170), 
	.A(n168));
   INVX1 U442 (.Y(n148), 
	.A(n147));
   INVX1 U443 (.Y(n130), 
	.A(n129));
   INVX1 U445 (.Y(n136), 
	.A(sboxw[25]));
   INVX1 U446 (.Y(n131), 
	.A(n128));
   INVX1 U447 (.Y(n162), 
	.A(n163));
   INVX1 U448 (.Y(n151), 
	.A(sboxw[16]));
   NOR2X1 U449 (.Y(n577), 
	.B(n130), 
	.A(n1583));
   NOR2X1 U450 (.Y(n931), 
	.B(n143), 
	.A(n211));
   NOR2X1 U451 (.Y(n348), 
	.B(n162), 
	.A(n1559));
   OAI32X1 U452 (.Y(n906), 
	.B1(n600), 
	.B0(n32), 
	.A2(n128), 
	.A1(n907), 
	.A0(n1583));
   AOI21X1 U453 (.Y(n907), 
	.B0(n40), 
	.A1(n11), 
	.A0(n730));
   NAND2X1 U454 (.Y(n631), 
	.B(n1583), 
	.A(n1593));
   NAND2X1 U455 (.Y(n985), 
	.B(n211), 
	.A(n56));
   NAND2X1 U456 (.Y(n402), 
	.B(n1559), 
	.A(n57));
   NOR3X1 U457 (.Y(n578), 
	.C(n4), 
	.B(n30), 
	.A(n604));
   AOI31X1 U458 (.Y(n875), 
	.B0(n581), 
	.A2(n66), 
	.A1(n129), 
	.A0(n138));
   AOI31X1 U459 (.Y(n1224), 
	.B0(n935), 
	.A2(n203), 
	.A1(n142), 
	.A0(n151));
   AOI31X1 U460 (.Y(n1129), 
	.B0(n352), 
	.A2(n1551), 
	.A1(n161), 
	.A0(n169));
   NAND2X1 U461 (.Y(n767), 
	.B(n1583), 
	.A(n1590));
   NAND2X1 U462 (.Y(n1088), 
	.B(n211), 
	.A(n204));
   NAND2X1 U463 (.Y(n505), 
	.B(n1559), 
	.A(n1552));
   NOR3XL U464 (.Y(n795), 
	.C(n4), 
	.B(n131), 
	.A(n662));
   NOR3XL U465 (.Y(n1144), 
	.C(n15), 
	.B(n143), 
	.A(n1016));
   NOR3XL U466 (.Y(n533), 
	.C(n16), 
	.B(sboxw[5]), 
	.A(n433));
   INVX1 U467 (.Y(n1587), 
	.A(n841));
   NAND2X1 U468 (.Y(n661), 
	.B(sboxw[24]), 
	.A(n67));
   NAND2X1 U469 (.Y(n1015), 
	.B(n150), 
	.A(n199));
   NAND2X1 U470 (.Y(n432), 
	.B(sboxw[0]), 
	.A(n1547));
   OAI211XL U471 (.Y(n710), 
	.C0(n573), 
	.B0(n611), 
	.A1(n4), 
	.A0(n576));
   NAND2X1 U472 (.Y(n600), 
	.B(n1578), 
	.A(n1590));
   NAND2X1 U473 (.Y(n595), 
	.B(n135), 
	.A(n66));
   NAND2X1 U474 (.Y(n582), 
	.B(n135), 
	.A(n1586));
   NAND3XL U475 (.Y(n287), 
	.C(n290), 
	.B(n1515), 
	.A(n25));
   INVX1 U476 (.Y(n216), 
	.A(n1435));
   NOR3X1 U477 (.Y(n1461), 
	.C(n60), 
	.B(n54), 
	.A(n318));
   NAND3X1 U478 (.Y(n846), 
	.C(n730), 
	.B(n1583), 
	.A(n122));
   NAND3X1 U479 (.Y(n1195), 
	.C(n1051), 
	.B(n211), 
	.A(n119));
   NAND3X1 U480 (.Y(n703), 
	.C(n468), 
	.B(n1559), 
	.A(n116));
   AOI21X1 U481 (.Y(n654), 
	.B0(n67), 
	.A1(n1593), 
	.A0(n136));
   AOI21X1 U482 (.Y(n1008), 
	.B0(n199), 
	.A1(n56), 
	.A0(n146));
   AOI21X1 U483 (.Y(n425), 
	.B0(n1547), 
	.A1(n57), 
	.A0(n167));
   NAND2X1 U484 (.Y(n734), 
	.B(n137), 
	.A(n63));
   NAND2X1 U485 (.Y(n472), 
	.B(sboxw[0]), 
	.A(n1536));
   NAND2X1 U486 (.Y(n594), 
	.B(n576), 
	.A(n67));
   NAND2X1 U487 (.Y(n948), 
	.B(n930), 
	.A(n199));
   NAND2X1 U488 (.Y(n365), 
	.B(n347), 
	.A(n1547));
   NAND3X1 U489 (.Y(n1414), 
	.C(n1102), 
	.B(n156), 
	.A(n1331));
   NAND2X1 U490 (.Y(n575), 
	.B(n1590), 
	.A(sboxw[24]));
   NAND2X1 U491 (.Y(n929), 
	.B(n204), 
	.A(n150));
   NAND2X1 U492 (.Y(n346), 
	.B(n1552), 
	.A(sboxw[0]));
   INVX1 U493 (.Y(n1595), 
	.A(n625));
   INVX1 U494 (.Y(n173), 
	.A(n979));
   INVX1 U495 (.Y(n1520), 
	.A(n396));
   NAND2X1 U496 (.Y(n597), 
	.B(n136), 
	.A(n63));
   NAND2X1 U497 (.Y(n951), 
	.B(n146), 
	.A(n64));
   NAND2X1 U498 (.Y(n368), 
	.B(n167), 
	.A(n1536));
   NAND2X1 U499 (.Y(n282), 
	.B(n1507), 
	.A(n49));
   NOR2X1 U500 (.Y(n891), 
	.B(n32), 
	.A(n48));
   XNOR2X1 U501 (.Y(n48), 
	.B(n137), 
	.A(n1583));
   INVX1 U502 (.Y(n645), 
	.A(n290));
   AOI22X1 U503 (.Y(n873), 
	.B1(n35), 
	.B0(n789), 
	.A1(n11), 
	.A0(n638));
   AOI22X1 U504 (.Y(n1222), 
	.B1(n36), 
	.B0(n1138), 
	.A1(n8), 
	.A0(n992));
   AOI22X1 U505 (.Y(n1127), 
	.B1(n37), 
	.B0(n527), 
	.A1(n7), 
	.A0(n409));
   NAND2X1 U506 (.Y(n611), 
	.B(n1590), 
	.A(n35));
   INVX1 U507 (.Y(n1572), 
	.A(n811));
   INVX1 U508 (.Y(n206), 
	.A(n1160));
   INVX1 U509 (.Y(n1554), 
	.A(n549));
   AOI22X1 U510 (.Y(n861), 
	.B1(n121), 
	.B0(n63), 
	.A1(n138), 
	.A0(n1590));
   AOI22X1 U511 (.Y(n1210), 
	.B1(n118), 
	.B0(n64), 
	.A1(n151), 
	.A0(n204));
   AOI22X1 U512 (.Y(n1115), 
	.B1(n115), 
	.B0(n1536), 
	.A1(n169), 
	.A0(n1552));
   NAND2X1 U513 (.Y(n601), 
	.B(n638), 
	.A(n135));
   NAND2X1 U514 (.Y(n955), 
	.B(n992), 
	.A(n147));
   NAND2X1 U515 (.Y(n372), 
	.B(n409), 
	.A(n166));
   NAND2X1 U516 (.Y(n837), 
	.B(n135), 
	.A(n801));
   NAND2X1 U517 (.Y(n655), 
	.B(n11), 
	.A(n801));
   NAND2X1 U518 (.Y(n1009), 
	.B(n8), 
	.A(n1150));
   NAND2X1 U519 (.Y(n426), 
	.B(n7), 
	.A(n539));
   INVX1 U520 (.Y(n571), 
	.A(n1297));
   INVX1 U521 (.Y(n1573), 
	.A(n836));
   INVX1 U522 (.Y(n124), 
	.A(n23));
   AND2X2 U525 (.Y(n49), 
	.B(sboxw[13]), 
	.A(n1515));
   INVX1 U526 (.Y(n318), 
	.A(n49));
   INVX1 U527 (.Y(n143), 
	.A(n142));
   INVX1 U528 (.Y(n215), 
	.A(n1442));
   NAND2X1 U529 (.Y(n651), 
	.B(n137), 
	.A(n1588));
   NAND2X1 U530 (.Y(n1005), 
	.B(n150), 
	.A(n205));
   NAND2X1 U531 (.Y(n422), 
	.B(n168), 
	.A(n1553));
   INVX1 U532 (.Y(n167), 
	.A(sboxw[1]));
   INVX1 U534 (.Y(n156), 
	.A(n153));
   OAI222XL U535 (.Y(n961), 
	.C1(n142), 
	.C0(n966), 
	.B1(n965), 
	.B0(n143), 
	.A1(n951), 
	.A0(n953));
   AND3X2 U536 (.Y(n966), 
	.C(n969), 
	.B(n968), 
	.A(n967));
   AOI222X1 U537 (.Y(n967), 
	.C1(n187), 
	.C0(n970), 
	.B1(n942), 
	.B0(n120), 
	.A1(n198), 
	.A0(n33));
   OAI221XL U538 (.Y(n1249), 
	.C0(n1250), 
	.B1(n1026), 
	.B0(n151), 
	.A1(n1163), 
	.A0(n33));
   AOI22X1 U539 (.Y(n1250), 
	.B1(n146), 
	.B0(n195), 
	.A1(n203), 
	.A0(n38));
   OAI221XL U540 (.Y(n1493), 
	.C0(n1494), 
	.B1(n443), 
	.B0(n170), 
	.A1(n552), 
	.A0(n34));
   AOI22X1 U541 (.Y(n1494), 
	.B1(n167), 
	.B0(n1543), 
	.A1(n1551), 
	.A0(n39));
   AOI222X1 U542 (.Y(n474), 
	.C1(n1526), 
	.C0(n31), 
	.B1(n160), 
	.B0(n476), 
	.A1(n475), 
	.A0(n159));
   OAI21XL U543 (.Y(n476), 
	.B0(n386), 
	.A1(n116), 
	.A0(n21));
   OAI211X1 U544 (.Y(n475), 
	.C0(n479), 
	.B0(n471), 
	.A1(n117), 
	.A0(n3));
   AOI22X1 U545 (.Y(n479), 
	.B1(n166), 
	.B0(n1536), 
	.A1(n117), 
	.A0(n1547));
   OAI221XL U546 (.Y(n824), 
	.C0(n826), 
	.B1(n781), 
	.B0(n135), 
	.A1(n583), 
	.A0(n576));
   OAI221XL U547 (.Y(n1173), 
	.C0(n1175), 
	.B1(n18), 
	.B0(n147), 
	.A1(n937), 
	.A0(n930));
   OAI221XL U548 (.Y(n681), 
	.C0(n683), 
	.B1(n19), 
	.B0(sboxw[1]), 
	.A1(n354), 
	.A0(n347));
   AOI222X1 U549 (.Y(n1057), 
	.C1(n179), 
	.C0(n29), 
	.B1(n142), 
	.B0(n1059), 
	.A1(n1058), 
	.A0(n143));
   OAI21XL U550 (.Y(n1059), 
	.B0(n969), 
	.A1(n119), 
	.A0(n20));
   OAI211X1 U551 (.Y(n1058), 
	.C0(n1062), 
	.B0(n1054), 
	.A1(n120), 
	.A0(n1));
   AOI22X1 U552 (.Y(n1062), 
	.B1(n147), 
	.B0(n64), 
	.A1(n120), 
	.A0(n199));
   OAI2BB2X1 U553 (.Y(n1170), 
	.B1(n1011), 
	.B0(n1171), 
	.A1N(n173), 
	.A0N(n1172));
   AOI211X1 U554 (.Y(n1171), 
	.C0(n1177), 
	.B0(n1176), 
	.A1(n148), 
	.A0(n198));
   NAND4BXL U555 (.Y(n1172), 
	.D(n1069), 
	.C(n1090), 
	.B(n1174), 
	.AN(n1173));
   OAI222XL U556 (.Y(n1176), 
	.C1(n120), 
	.C0(n20), 
	.B1(n1163), 
	.B0(n27), 
	.A1(n1026), 
	.A0(n930));
   OAI2BB2X1 U557 (.Y(n821), 
	.B1(n657), 
	.B0(n822), 
	.A1N(n1595), 
	.A0N(n823));
   AOI211X1 U558 (.Y(n822), 
	.C0(n828), 
	.B0(n827), 
	.A1(n136), 
	.A0(n1574));
   NAND4BXL U559 (.Y(n823), 
	.D(n748), 
	.C(n769), 
	.B(n825), 
	.AN(n824));
   OAI222XL U560 (.Y(n827), 
	.C1(n123), 
	.C0(n2), 
	.B1(n814), 
	.B0(n26), 
	.A1(n14), 
	.A0(n576));
   OAI2BB2X1 U561 (.Y(n678), 
	.B1(n428), 
	.B0(n679), 
	.A1N(n1520), 
	.A0N(n680));
   AOI211X1 U562 (.Y(n679), 
	.C0(n685), 
	.B0(n684), 
	.A1(n167), 
	.A0(n1546));
   NAND4BXL U563 (.Y(n680), 
	.D(n486), 
	.C(n507), 
	.B(n682), 
	.AN(n681));
   OAI222XL U564 (.Y(n684), 
	.C1(n117), 
	.C0(n21), 
	.B1(n552), 
	.B0(n28), 
	.A1(n443), 
	.A0(n347));
   OAI21XL U565 (.Y(n1245), 
	.B0(n1247), 
	.A1(n142), 
	.A0(n1246));
   AOI31X1 U566 (.Y(n1247), 
	.B0(n180), 
	.A2(n36), 
	.A1(n207), 
	.A0(n181));
   NOR4BX1 U567 (.Y(n1246), 
	.D(n960), 
	.C(n198), 
	.B(n1249), 
	.AN(n1248));
   AOI21X1 U568 (.Y(n1248), 
	.B0(n981), 
	.A1(n202), 
	.A0(n119));
   OAI21XL U569 (.Y(n1489), 
	.B0(n1491), 
	.A1(n161), 
	.A0(n1490));
   AOI31X1 U570 (.Y(n1491), 
	.B0(n1527), 
	.A2(n37), 
	.A1(n1555), 
	.A0(n1528));
   NOR4BX1 U571 (.Y(n1490), 
	.D(n377), 
	.C(n1546), 
	.B(n1493), 
	.AN(n1492));
   AOI21X1 U572 (.Y(n1492), 
	.B0(n398), 
	.A1(n1550), 
	.A0(n116));
   INVX1 U574 (.Y(n1585), 
	.A(n643));
   INVX1 U576 (.Y(n195), 
	.A(n997));
   INVX1 U578 (.Y(n1543), 
	.A(n414));
   NOR2X1 U579 (.Y(n1160), 
	.B(n1093), 
	.A(n1079));
   NOR2X1 U580 (.Y(n549), 
	.B(n510), 
	.A(n496));
   NOR2X1 U581 (.Y(n227), 
	.B(n243), 
	.A(n1342));
   AOI222XL U582 (.Y(n289), 
	.C1(n247), 
	.C0(n59), 
	.B1(n1503), 
	.B0(n50), 
	.A1(n23), 
	.A0(n1506));
   AOI222X1 U583 (.Y(n810), 
	.C1(n616), 
	.C0(n1575), 
	.B1(n139), 
	.B0(n780), 
	.A1(n1572), 
	.A0(n32));
   AOI222X1 U584 (.Y(n1159), 
	.C1(n970), 
	.C0(n190), 
	.B1(n151), 
	.B0(n1101), 
	.A1(n206), 
	.A0(n33));
   AOI222X1 U585 (.Y(n548), 
	.C1(n387), 
	.C0(n1538), 
	.B1(n169), 
	.B0(n518), 
	.A1(n1554), 
	.A0(n34));
   OAI222XL U586 (.Y(n1373), 
	.C1(n156), 
	.C0(n1376), 
	.B1(n1375), 
	.B0(n153), 
	.A1(n1265), 
	.A0(n24));
   AOI21X1 U587 (.Y(n1375), 
	.B0(n1302), 
	.A1(n60), 
	.A0(n50));
   AOI211X1 U588 (.Y(n1376), 
	.C0(n925), 
	.B0(n1377), 
	.A1(n1502), 
	.A0(n65));
   OAI22X1 U589 (.Y(n1377), 
	.B1(n17), 
	.B0(n65), 
	.A1(n1516), 
	.A0(n243));
   OAI222XL U590 (.Y(n1262), 
	.C1(n1265), 
	.C0(n240), 
	.B1(n1264), 
	.B0(n153), 
	.A1(sboxw[13]), 
	.A0(n1263));
   AOI221XL U591 (.Y(n1263), 
	.C0(n1266), 
	.B1(n24), 
	.B0(n58), 
	.A1(n1507), 
	.A0(n124));
   AOI211X1 U592 (.Y(n1264), 
	.C0(n1504), 
	.B0(n1501), 
	.A1(n1061), 
	.A0(n55));
   INVX1 U593 (.Y(n1504), 
	.A(n258));
   OAI32X1 U594 (.Y(n321), 
	.B1(n323), 
	.B0(n55), 
	.A2(n156), 
	.A1(n322), 
	.A0(n1515));
   AOI21XL U595 (.Y(n322), 
	.B0(n50), 
	.A1(n23), 
	.A0(n290));
   NOR2X1 U596 (.Y(n274), 
	.B(n230), 
	.A(n1342));
   NAND4X1 U597 (.Y(n700), 
	.D(n704), 
	.C(n703), 
	.B(n414), 
	.A(n1548));
   AOI221X1 U598 (.Y(n704), 
	.C0(n705), 
	.B1(n34), 
	.B0(n518), 
	.A1(n28), 
	.A0(n1546));
   AOI21X1 U599 (.Y(n705), 
	.B0(n167), 
	.A1(n431), 
	.A0(n16));
   OAI222XL U600 (.Y(n639), 
	.C1(n22), 
	.C0(n644), 
	.B1(n123), 
	.B0(n643), 
	.A1(n10), 
	.A0(n642));
   OAI222XL U601 (.Y(n993), 
	.C1(n999), 
	.C0(n998), 
	.B1(n120), 
	.B0(n997), 
	.A1(n6), 
	.A0(n996));
   OAI222XL U602 (.Y(n410), 
	.C1(n416), 
	.C0(n415), 
	.B1(n117), 
	.B0(n414), 
	.A1(n5), 
	.A0(n9));
   NAND4BXL U603 (.Y(n1030), 
	.D(n1033), 
	.C(n200), 
	.B(n959), 
	.AN(n943));
   AOI211X1 U604 (.Y(n1033), 
	.C0(n1034), 
	.B0(n210), 
	.A1(n29), 
	.A0(n187));
   AOI21X1 U605 (.Y(n1034), 
	.B0(n118), 
	.A1(n985), 
	.A0(n1026));
   INVX1 U606 (.Y(n210), 
	.A(n1035));
   NAND4X1 U607 (.Y(n1356), 
	.D(n1358), 
	.C(n1357), 
	.B(n248), 
	.A(n259));
   AOI21X1 U608 (.Y(n1357), 
	.B0(n273), 
	.A1(n1365), 
	.A0(n49));
   AOI211XL U609 (.Y(n1358), 
	.C0(n1360), 
	.B0(n1359), 
	.A1(n23), 
	.A0(n739));
   OAI21XL U610 (.Y(n1365), 
	.B0(n24), 
	.A1(n1511), 
	.A0(n55));
   AOI221XL U611 (.Y(n1419), 
	.C0(n989), 
	.B1(n247), 
	.B0(n1277), 
	.A1(n23), 
	.A0(n635));
   INVX1 U612 (.Y(n989), 
	.A(n259));
   OAI222XL U613 (.Y(n1293), 
	.C1(sboxw[13]), 
	.C0(n1299), 
	.B1(n1298), 
	.B0(n153), 
	.A1(n1297), 
	.A0(n318));
   NOR3BX1 U614 (.Y(n1299), 
	.C(n1302), 
	.B(n1301), 
	.AN(n1300));
   OAI222XL U615 (.Y(n378), 
	.C1(n161), 
	.C0(n383), 
	.B1(n382), 
	.B0(n162), 
	.A1(n368), 
	.A0(n370));
   AND3X2 U616 (.Y(n383), 
	.C(n386), 
	.B(n385), 
	.A(n384));
   AOI222X1 U617 (.Y(n384), 
	.C1(n1534), 
	.C0(n387), 
	.B1(n359), 
	.B0(n117), 
	.A1(n1546), 
	.A0(n34));
   OAI222XL U618 (.Y(n812), 
	.C1(n576), 
	.C0(n740), 
	.B1(n138), 
	.B0(n814), 
	.A1(n644), 
	.A0(n22));
   OAI222XL U619 (.Y(n1161), 
	.C1(n930), 
	.C0(n1), 
	.B1(n151), 
	.B0(n1163), 
	.A1(n998), 
	.A0(n999));
   OAI222XL U620 (.Y(n550), 
	.C1(n347), 
	.C0(n3), 
	.B1(n169), 
	.B0(n552), 
	.A1(n415), 
	.A0(n416));
   OAI221XL U621 (.Y(n900), 
	.C0(n901), 
	.B1(n14), 
	.B0(n138), 
	.A1(n814), 
	.A0(n32));
   AOI22X1 U622 (.Y(n901), 
	.B1(n136), 
	.B0(n1585), 
	.A1(n66), 
	.A0(n40));
   NOR2X1 U623 (.Y(n960), 
	.B(n18), 
	.A(n8));
   NOR2X1 U624 (.Y(n377), 
	.B(n19), 
	.A(n7));
   AOI222X1 U625 (.Y(n294), 
	.C1(n1516), 
	.C0(n273), 
	.B1(n156), 
	.B0(n296), 
	.A1(n295), 
	.A0(n153));
   OAI221XL U626 (.Y(n296), 
	.C0(n298), 
	.B1(n25), 
	.B0(n13), 
	.A1(n243), 
	.A0(n297));
   NAND4X1 U627 (.Y(n295), 
	.D(n300), 
	.C(n299), 
	.B(n246), 
	.A(n248));
   AOI21X1 U628 (.Y(n299), 
	.B0(n303), 
	.A1(n290), 
	.A0(n302));
   NOR2X1 U629 (.Y(n1266), 
	.B(n54), 
	.A(n12));
   NOR2X1 U630 (.Y(n589), 
	.B(n35), 
	.A(n740));
   NOR2X1 U631 (.Y(n943), 
	.B(n36), 
	.A(n1));
   NOR2X1 U632 (.Y(n360), 
	.B(n37), 
	.A(n3));
   NOR2X1 U633 (.Y(n1150), 
	.B(n20), 
	.A(n953));
   NOR2X1 U634 (.Y(n539), 
	.B(n21), 
	.A(n370));
   OAI221XL U635 (.Y(n894), 
	.C0(n904), 
	.B1(n814), 
	.B0(n616), 
	.A1(n903), 
	.A0(n130));
   AOI21X1 U636 (.Y(n904), 
	.B0(n906), 
	.A1(n905), 
	.A0(n1581));
   AOI221X1 U637 (.Y(n903), 
	.C0(n778), 
	.B1(n122), 
	.B0(n1586), 
	.A1(n121), 
	.A0(n1585));
   OAI221XL U638 (.Y(n905), 
	.C0(n734), 
	.B1(n4), 
	.B0(sboxw[24]), 
	.A1(n576), 
	.A0(n2));
   OAI221XL U639 (.Y(n1243), 
	.C0(n1253), 
	.B1(n1163), 
	.B0(n970), 
	.A1(n1252), 
	.A0(n143));
   AOI21X1 U640 (.Y(n1253), 
	.B0(n1255), 
	.A1(n1254), 
	.A0(n181));
   AOI221X1 U641 (.Y(n1252), 
	.C0(n1099), 
	.B1(n6), 
	.B0(n61), 
	.A1(n118), 
	.A0(n195));
   OAI221XL U642 (.Y(n1254), 
	.C0(n1055), 
	.B1(n15), 
	.B0(sboxw[16]), 
	.A1(n930), 
	.A0(n20));
   OAI221XL U643 (.Y(n1487), 
	.C0(n1497), 
	.B1(n552), 
	.B0(n387), 
	.A1(n1496), 
	.A0(n159));
   AOI21X1 U644 (.Y(n1497), 
	.B0(n1499), 
	.A1(n1498), 
	.A0(n1528));
   AOI221X1 U645 (.Y(n1496), 
	.C0(n516), 
	.B1(n5), 
	.B0(n62), 
	.A1(n115), 
	.A0(n1543));
   OAI221XL U646 (.Y(n1498), 
	.C0(n472), 
	.B1(n16), 
	.B0(sboxw[0]), 
	.A1(n347), 
	.A0(n21));
   OAI221XL U647 (.Y(n1305), 
	.C0(n1317), 
	.B1(n1316), 
	.B0(n153), 
	.A1(n156), 
	.A0(n1315));
   AOI22X1 U648 (.Y(n1317), 
	.B1(n65), 
	.B0(n227), 
	.A1(n50), 
	.A0(n274));
   AOI211X1 U649 (.Y(n1315), 
	.C0(n1501), 
	.B0(n1322), 
	.A1(n1516), 
	.A0(n1102));
   AOI211X1 U650 (.Y(n1316), 
	.C0(n1319), 
	.B0(n1318), 
	.A1(n1495), 
	.A0(n127));
   OAI221XL U651 (.Y(n305), 
	.C0(n320), 
	.B1(n319), 
	.B0(n153), 
	.A1(n318), 
	.A0(n317));
   AOI221X1 U652 (.Y(n317), 
	.C0(n519), 
	.B1(n240), 
	.B0(n60), 
	.A1(n1517), 
	.A0(n1102));
   AOI221XL U653 (.Y(n319), 
	.C0(n232), 
	.B1(n25), 
	.B0(n59), 
	.A1(n23), 
	.A0(n1061));
   AOI21X1 U654 (.Y(n320), 
	.B0(n321), 
	.A1(n227), 
	.A0(n55));
   OAI221XL U655 (.Y(n306), 
	.C0(n316), 
	.B1(n243), 
	.B0(n297), 
	.A1(n247), 
	.A0(n12));
   OAI221XL U656 (.Y(n619), 
	.C0(n637), 
	.B1(n636), 
	.B0(sboxw[29]), 
	.A1(n128), 
	.A0(n1563));
   AOI22X1 U657 (.Y(n637), 
	.B1(n638), 
	.B0(n40), 
	.A1(n30), 
	.A0(n1577));
   INVX1 U658 (.Y(n1563), 
	.A(n646));
   AOI211X1 U659 (.Y(n636), 
	.C0(n640), 
	.B0(n639), 
	.A1(n576), 
	.A0(n1576));
   OAI221XL U660 (.Y(n390), 
	.C0(n408), 
	.B1(n407), 
	.B0(sboxw[5]), 
	.A1(n160), 
	.A0(n1535));
   AOI22X1 U661 (.Y(n408), 
	.B1(n409), 
	.B0(n39), 
	.A1(n31), 
	.A0(n1531));
   INVX1 U662 (.Y(n1535), 
	.A(n417));
   AOI211X1 U663 (.Y(n407), 
	.C0(n411), 
	.B0(n410), 
	.A1(n347), 
	.A0(n1550));
   OAI221XL U664 (.Y(n310), 
	.C0(n315), 
	.B1(n254), 
	.B0(n1517), 
	.A1(n314), 
	.A0(n55));
   AOI211X1 U665 (.Y(n852), 
	.C0(n858), 
	.B0(n857), 
	.A1(n856), 
	.A0(n1578));
   OAI221XL U666 (.Y(n856), 
	.C0(n861), 
	.B1(n139), 
	.B0(n22), 
	.A1(n4), 
	.A0(n40));
   AOI31X1 U667 (.Y(n857), 
	.B0(n130), 
	.A2(n860), 
	.A1(n654), 
	.A0(n859));
   AOI31X1 U668 (.Y(n858), 
	.B0(n128), 
	.A2(n596), 
	.A1(n769), 
	.A0(n718));
   AOI211X1 U669 (.Y(n1201), 
	.C0(n1207), 
	.B0(n1206), 
	.A1(n1205), 
	.A0(n185));
   OAI221XL U670 (.Y(n1205), 
	.C0(n1210), 
	.B1(n151), 
	.B0(n999), 
	.A1(n15), 
	.A0(n38));
   AOI31X1 U671 (.Y(n1206), 
	.B0(sboxw[21]), 
	.A2(n1209), 
	.A1(n1008), 
	.A0(n1208));
   AOI31X1 U672 (.Y(n1207), 
	.B0(n142), 
	.A2(n950), 
	.A1(n1090), 
	.A0(n1039));
   AOI211X1 U673 (.Y(n1106), 
	.C0(n1112), 
	.B0(n1111), 
	.A1(n1110), 
	.A0(n1532));
   OAI221XL U674 (.Y(n1110), 
	.C0(n1115), 
	.B1(n169), 
	.B0(n416), 
	.A1(n16), 
	.A0(n39));
   AOI31X1 U675 (.Y(n1111), 
	.B0(sboxw[5]), 
	.A2(n1114), 
	.A1(n425), 
	.A0(n1113));
   AOI31X1 U676 (.Y(n1112), 
	.B0(n160), 
	.A2(n367), 
	.A1(n507), 
	.A0(n456));
   OAI221XL U677 (.Y(n973), 
	.C0(n991), 
	.B1(n990), 
	.B0(sboxw[21]), 
	.A1(n142), 
	.A0(n188));
   AOI22X1 U678 (.Y(n991), 
	.B1(n992), 
	.B0(n38), 
	.A1(n29), 
	.A0(n184));
   INVX1 U679 (.Y(n188), 
	.A(n1000));
   AOI211X1 U680 (.Y(n990), 
	.C0(n994), 
	.B0(n993), 
	.A1(n930), 
	.A0(n202));
   AOI211X1 U681 (.Y(n851), 
	.C0(n863), 
	.B0(n862), 
	.A1(n35), 
	.A0(n1574));
   OAI222XL U682 (.Y(n862), 
	.C1(n123), 
	.C0(n642), 
	.B1(n14), 
	.B0(sboxw[24]), 
	.A1(n740), 
	.A0(n40));
   OAI21XL U683 (.Y(n863), 
	.B0(n864), 
	.A1(n829), 
	.A0(n26));
   OAI21XL U684 (.Y(n864), 
	.B0(n137), 
	.A1(n1585), 
	.A0(n1576));
   AOI211X1 U685 (.Y(n1200), 
	.C0(n1212), 
	.B0(n1211), 
	.A1(n36), 
	.A0(n198));
   OAI222XL U686 (.Y(n1211), 
	.C1(n120), 
	.C0(n996), 
	.B1(n1026), 
	.B0(sboxw[16]), 
	.A1(n1), 
	.A0(n38));
   OAI21XL U687 (.Y(n1212), 
	.B0(n1213), 
	.A1(n1178), 
	.A0(n27));
   OAI21XL U688 (.Y(n1213), 
	.B0(n150), 
	.A1(n195), 
	.A0(n202));
   AOI211X1 U689 (.Y(n1105), 
	.C0(n1117), 
	.B0(n1116), 
	.A1(n37), 
	.A0(n1546));
   OAI222XL U690 (.Y(n1116), 
	.C1(n117), 
	.C0(n9), 
	.B1(n443), 
	.B0(sboxw[0]), 
	.A1(n3), 
	.A0(n39));
   OAI21XL U691 (.Y(n1117), 
	.B0(n1118), 
	.A1(n686), 
	.A0(n28));
   OAI21XL U692 (.Y(n1118), 
	.B0(n168), 
	.A1(n1543), 
	.A0(n1550));
   NOR2BX1 U693 (.Y(n286), 
	.B(n153), 
	.AN(n1314));
   NOR2X1 U694 (.Y(n263), 
	.B(n1374), 
	.A(n1516));
   NOR2XL U695 (.Y(n1341), 
	.B(n1374), 
	.A(n23));
   NOR2X1 U696 (.Y(n1364), 
	.B(n12), 
	.A(n125));
   NOR2X1 U697 (.Y(n725), 
	.B(n26), 
	.A(n740));
   NOR2X1 U698 (.Y(n1046), 
	.B(n27), 
	.A(n1));
   NOR2X1 U699 (.Y(n463), 
	.B(n28), 
	.A(n3));
   AOI222X1 U700 (.Y(n736), 
	.C1(n1579), 
	.C0(n30), 
	.B1(n128), 
	.B0(n738), 
	.A1(n737), 
	.A0(n130));
   OAI21XL U701 (.Y(n738), 
	.B0(n615), 
	.A1(n122), 
	.A0(n2));
   OAI211X1 U702 (.Y(n737), 
	.C0(n741), 
	.B0(n733), 
	.A1(n123), 
	.A0(n740));
   AOI22X1 U703 (.Y(n741), 
	.B1(n135), 
	.B0(n63), 
	.A1(n123), 
	.A0(n67));
   OAI211X1 U704 (.Y(n834), 
	.C0(n839), 
	.B0(n614), 
	.A1(n14), 
	.A0(n576));
   AOI211X1 U705 (.Y(n839), 
	.C0(n840), 
	.B0(n668), 
	.A1(n616), 
	.A0(n1576));
   NOR3X1 U706 (.Y(n840), 
	.C(n811), 
	.B(n30), 
	.A(n1594));
   OAI211X1 U707 (.Y(n1183), 
	.C0(n1188), 
	.B0(n968), 
	.A1(n1026), 
	.A0(n930));
   AOI211X1 U708 (.Y(n1188), 
	.C0(n1189), 
	.B0(n1022), 
	.A1(n970), 
	.A0(n202));
   NOR3X1 U709 (.Y(n1189), 
	.C(n1160), 
	.B(n29), 
	.A(n197));
   OAI211X1 U710 (.Y(n691), 
	.C0(n696), 
	.B0(n385), 
	.A1(n443), 
	.A0(n347));
   AOI211X1 U711 (.Y(n696), 
	.C0(n697), 
	.B0(n439), 
	.A1(n387), 
	.A0(n1550));
   NOR3X1 U712 (.Y(n697), 
	.C(n549), 
	.B(n31), 
	.A(n1545));
   OAI211X1 U713 (.Y(n842), 
	.C0(n826), 
	.B0(n661), 
	.A1(n740), 
	.A0(sboxw[25]));
   OAI211X1 U714 (.Y(n1191), 
	.C0(n1175), 
	.B0(n1015), 
	.A1(n1), 
	.A0(n147));
   OAI211X1 U715 (.Y(n699), 
	.C0(n683), 
	.B0(n432), 
	.A1(n3), 
	.A0(sboxw[1]));
   OAI211X1 U716 (.Y(n1239), 
	.C0(n949), 
	.B0(n959), 
	.A1(n996), 
	.A0(n1240));
   OAI211X1 U717 (.Y(n1483), 
	.C0(n366), 
	.B0(n376), 
	.A1(n9), 
	.A0(n1484));
   NAND2X1 U718 (.Y(n1278), 
	.B(n1394), 
	.A(n314));
   INVX1 U719 (.Y(n1502), 
	.A(n12));
   NOR4BX1 U720 (.Y(n755), 
	.D(n1588), 
	.C(n757), 
	.B(n627), 
	.AN(n756));
   AOI2BB1X1 U721 (.Y(n757), 
	.B0(n30), 
	.A1N(n629), 
	.A0N(n1593));
   AOI222X1 U722 (.Y(n756), 
	.C1(n40), 
	.C0(n1590), 
	.B1(n758), 
	.B0(n35), 
	.A1(n1582), 
	.A0(n137));
   NOR4BX1 U723 (.Y(n1076), 
	.D(n205), 
	.C(n1078), 
	.B(n981), 
	.AN(n1077));
   AOI2BB1X1 U724 (.Y(n1078), 
	.B0(n29), 
	.A1N(n983), 
	.A0N(n56));
   AOI222X1 U725 (.Y(n1077), 
	.C1(n38), 
	.C0(n204), 
	.B1(n1079), 
	.B0(n36), 
	.A1(n187), 
	.A0(sboxw[16]));
   NOR4BX1 U726 (.Y(n493), 
	.D(n1553), 
	.C(n495), 
	.B(n398), 
	.AN(n494));
   AOI2BB1X1 U727 (.Y(n495), 
	.B0(n31), 
	.A1N(n400), 
	.A0N(n57));
   AOI222X1 U728 (.Y(n494), 
	.C1(n39), 
	.C0(n1552), 
	.B1(n496), 
	.B0(n37), 
	.A1(n1534), 
	.A0(n168));
   AOI31XL U729 (.Y(n1360), 
	.B0(n1342), 
	.A2(n1298), 
	.A1(n243), 
	.A0(n1361));
   NOR4X1 U730 (.Y(n1391), 
	.D(n313), 
	.C(n1393), 
	.B(n1392), 
	.A(n1508));
   AOI2BB1X1 U731 (.Y(n1393), 
	.B0(n65), 
	.A1N(n1313), 
	.A0N(n1507));
   AOI31X1 U732 (.Y(n1043), 
	.B0(n958), 
	.A2(n965), 
	.A1(n996), 
	.A0(n1023));
   AOI31X1 U733 (.Y(n460), 
	.B0(n375), 
	.A2(n382), 
	.A1(n9), 
	.A0(n440));
   OAI21XL U734 (.Y(n1301), 
	.B0(n1284), 
	.A1(n246), 
	.A0(n50));
   AOI22X1 U735 (.Y(n315), 
	.B1(n1061), 
	.B0(n1516), 
	.A1(n54), 
	.A0(n1507));
   AOI31X1 U736 (.Y(n1441), 
	.B0(n1364), 
	.A2(n1510), 
	.A1(n1251), 
	.A0(n55));
   AOI31X1 U737 (.Y(n1164), 
	.B0(n1046), 
	.A2(n1160), 
	.A1(n197), 
	.A0(n33));
   AOI31X1 U738 (.Y(n553), 
	.B0(n463), 
	.A2(n549), 
	.A1(n1545), 
	.A0(n34));
   AOI31X1 U739 (.Y(n803), 
	.B0(n625), 
	.A2(n806), 
	.A1(n805), 
	.A0(n804));
   AOI222X1 U740 (.Y(n806), 
	.C1(n67), 
	.C0(n40), 
	.B1(n139), 
	.B0(n1586), 
	.A1(n1590), 
	.A0(n663));
   AOI22X1 U741 (.Y(n804), 
	.B1(n30), 
	.B0(n1582), 
	.A1(n137), 
	.A0(n1575));
   AOI21X1 U742 (.Y(n805), 
	.B0(n1565), 
	.A1(n576), 
	.A0(n1574));
   AOI31X1 U743 (.Y(n1152), 
	.B0(n979), 
	.A2(n1155), 
	.A1(n1154), 
	.A0(n1153));
   AOI222X1 U744 (.Y(n1155), 
	.C1(n199), 
	.C0(n38), 
	.B1(n151), 
	.B0(n61), 
	.A1(n204), 
	.A0(n1017));
   AOI22X1 U745 (.Y(n1153), 
	.B1(n29), 
	.B0(n187), 
	.A1(n150), 
	.A0(n190));
   AOI21X1 U746 (.Y(n1154), 
	.B0(n194), 
	.A1(n930), 
	.A0(n198));
   AOI31X1 U747 (.Y(n541), 
	.B0(n396), 
	.A2(n544), 
	.A1(n543), 
	.A0(n542));
   AOI222X1 U748 (.Y(n544), 
	.C1(n1547), 
	.C0(n39), 
	.B1(n170), 
	.B0(n62), 
	.A1(n1552), 
	.A0(n434));
   AOI22X1 U749 (.Y(n542), 
	.B1(n31), 
	.B0(n1534), 
	.A1(n168), 
	.A0(n1538));
   AOI21X1 U750 (.Y(n543), 
	.B0(n1542), 
	.A1(n347), 
	.A0(n1546));
   AOI31X1 U751 (.Y(n650), 
	.B0(n565), 
	.A2(n1561), 
	.A1(n652), 
	.A0(n651));
   INVX1 U752 (.Y(n1561), 
	.A(n653));
   OAI21XL U753 (.Y(n653), 
	.B0(n654), 
	.A1(n644), 
	.A0(n642));
   AOI31X1 U754 (.Y(n1004), 
	.B0(n919), 
	.A2(n189), 
	.A1(n1006), 
	.A0(n1005));
   INVX1 U755 (.Y(n189), 
	.A(n1007));
   OAI21XL U756 (.Y(n1007), 
	.B0(n1008), 
	.A1(n998), 
	.A0(n996));
   AOI31X1 U757 (.Y(n421), 
	.B0(n336), 
	.A2(n1537), 
	.A1(n423), 
	.A0(n422));
   INVX1 U758 (.Y(n1537), 
	.A(n424));
   OAI21XL U759 (.Y(n424), 
	.B0(n425), 
	.A1(n415), 
	.A0(n9));
   NAND2XL U760 (.Y(n259), 
	.B(n24), 
	.A(n1061));
   NAND2X1 U761 (.Y(n252), 
	.B(n1290), 
	.A(n17));
   NOR2X1 U762 (.Y(n1190), 
	.B(n150), 
	.A(n18));
   NOR2X1 U763 (.Y(n698), 
	.B(sboxw[0]), 
	.A(n19));
   NOR2X1 U764 (.Y(n1016), 
	.B(n38), 
	.A(n988));
   NOR2X1 U765 (.Y(n433), 
	.B(n39), 
	.A(n405));
   NOR2X1 U766 (.Y(n271), 
	.B(n153), 
	.A(n254));
   NOR2X1 U767 (.Y(n935), 
	.B(n143), 
	.A(n1026));
   NOR2X1 U768 (.Y(n352), 
	.B(sboxw[5]), 
	.A(n443));
   OAI22X1 U769 (.Y(n1359), 
	.B1(n1363), 
	.B0(n153), 
	.A1(sboxw[13]), 
	.A0(n1362));
   AOI21X1 U770 (.Y(n1362), 
	.B0(n1506), 
	.A1(n1517), 
	.A0(n1313));
   AOI21XL U771 (.Y(n1363), 
	.B0(n1364), 
	.A1(n247), 
	.A0(n58));
   AOI22XL U772 (.Y(n269), 
	.B1(n25), 
	.B0(n406), 
	.A1(n272), 
	.A0(n153));
   OAI22X1 U773 (.Y(n272), 
	.B1(n12), 
	.B0(n1517), 
	.A1(n17), 
	.A0(n65));
   AOI22XL U774 (.Y(n236), 
	.B1(n23), 
	.B0(n1061), 
	.A1(n125), 
	.A0(n635));
   OAI21XL U775 (.Y(n1421), 
	.B0(n153), 
	.A1(n1425), 
	.A0(n1424));
   OAI222XL U776 (.Y(n1425), 
	.C1(n1514), 
	.C0(n242), 
	.B1(n24), 
	.B0(n254), 
	.A1(n17), 
	.A0(n50));
   OAI222XL U777 (.Y(n1424), 
	.C1(n1290), 
	.C0(n1516), 
	.B1(n240), 
	.B0(n1426), 
	.A1(n262), 
	.A0(n23));
   INVX1 U778 (.Y(n1514), 
	.A(n1321));
   NAND2X1 U779 (.Y(n1277), 
	.B(n1311), 
	.A(n254));
   NAND2X1 U780 (.Y(n920), 
	.B(n1088), 
	.A(n1026));
   NAND2X1 U781 (.Y(n337), 
	.B(n505), 
	.A(n443));
   NAND4X1 U782 (.Y(n889), 
	.D(n893), 
	.C(n892), 
	.B(n643), 
	.A(n718));
   AOI21X1 U783 (.Y(n892), 
	.B0(n1571), 
	.A1(n730), 
	.A0(n634));
   AOI222X1 U784 (.Y(n893), 
	.C1(n30), 
	.C0(n1574), 
	.B1(n35), 
	.B0(n780), 
	.A1(n137), 
	.A0(n1591));
   INVX1 U785 (.Y(n1571), 
	.A(n830));
   NAND4X1 U786 (.Y(n1238), 
	.D(n1242), 
	.C(n1241), 
	.B(n997), 
	.A(n1039));
   AOI21X1 U787 (.Y(n1241), 
	.B0(n208), 
	.A1(n1051), 
	.A0(n988));
   AOI222X1 U788 (.Y(n1242), 
	.C1(n29), 
	.C0(n198), 
	.B1(n36), 
	.B0(n1101), 
	.A1(n150), 
	.A0(n196));
   INVX1 U789 (.Y(n208), 
	.A(n1179));
   NAND4X1 U790 (.Y(n1482), 
	.D(n1486), 
	.C(n1485), 
	.B(n414), 
	.A(n456));
   AOI21X1 U791 (.Y(n1485), 
	.B0(n1556), 
	.A1(n468), 
	.A0(n405));
   AOI222X1 U792 (.Y(n1486), 
	.C1(n31), 
	.C0(n1546), 
	.B1(n37), 
	.B0(n518), 
	.A1(n168), 
	.A0(n1544));
   INVX1 U793 (.Y(n1556), 
	.A(n687));
   AOI21XL U794 (.Y(n288), 
	.B0(n1060), 
	.A1(n24), 
	.A0(n739));
   NAND4X1 U795 (.Y(n1192), 
	.D(n1196), 
	.C(n1195), 
	.B(n997), 
	.A(n200));
   AOI221X1 U796 (.Y(n1196), 
	.C0(n1197), 
	.B1(n33), 
	.B0(n1101), 
	.A1(n27), 
	.A0(n198));
   AOI21X1 U797 (.Y(n1197), 
	.B0(n148), 
	.A1(n1014), 
	.A0(n15));
   NAND2X1 U798 (.Y(n1035), 
	.B(n33), 
	.A(n942));
   NAND2X1 U799 (.Y(n452), 
	.B(n34), 
	.A(n359));
   OAI21XL U800 (.Y(n1370), 
	.B0(n1371), 
	.A1(n1290), 
	.A0(n1516));
   NAND4X1 U801 (.Y(n1466), 
	.D(n1468), 
	.C(n287), 
	.B(n246), 
	.A(n1284));
   AOI221X1 U802 (.Y(n1468), 
	.C0(n1469), 
	.B1(n55), 
	.B0(n301), 
	.A1(n240), 
	.A0(n1503));
   AOI21X1 U803 (.Y(n1469), 
	.B0(n1516), 
	.A1(n1333), 
	.A0(n13));
   INVX1 U804 (.Y(n1564), 
	.A(n807));
   AOI22X1 U805 (.Y(n807), 
	.B1(n809), 
	.B0(n1596), 
	.A1(n808), 
	.A0(n1597));
   NAND4BXL U806 (.Y(n808), 
	.D(n813), 
	.C(n748), 
	.B(n596), 
	.AN(n812));
   NAND4X1 U807 (.Y(n809), 
	.D(n810), 
	.C(n651), 
	.B(n22), 
	.A(n768));
   INVX1 U808 (.Y(n1522), 
	.A(n545));
   AOI22X1 U809 (.Y(n545), 
	.B1(n547), 
	.B0(n1523), 
	.A1(n546), 
	.A0(n1524));
   NAND4BXL U810 (.Y(n546), 
	.D(n551), 
	.C(n486), 
	.B(n367), 
	.AN(n550));
   NAND4X1 U811 (.Y(n547), 
	.D(n548), 
	.C(n422), 
	.B(n416), 
	.A(n506));
   NAND4X1 U812 (.Y(n1307), 
	.D(n1310), 
	.C(n1309), 
	.B(n1308), 
	.A(n1289));
   AOI22X1 U813 (.Y(n1309), 
	.B1(n50), 
	.B0(n739), 
	.A1(n13), 
	.A0(n302));
   AOI222X1 U814 (.Y(n1310), 
	.C1(n1061), 
	.C0(n127), 
	.B1(n240), 
	.B0(n1502), 
	.A1(n1516), 
	.A0(n1507));
   NAND2X1 U815 (.Y(n1185), 
	.B(n142), 
	.A(n980));
   NAND2X1 U816 (.Y(n693), 
	.B(n161), 
	.A(n397));
   INVX1 U817 (.Y(n1568), 
	.A(n669));
   INVX1 U818 (.Y(n209), 
	.A(n1023));
   INVX1 U819 (.Y(n1557), 
	.A(n440));
   NAND4X1 U820 (.Y(n716), 
	.D(n720), 
	.C(n719), 
	.B(n718), 
	.A(n717));
   AOI21X1 U821 (.Y(n719), 
	.B0(n1579), 
	.A1(n726), 
	.A0(n1581));
   AOI211X1 U822 (.Y(n720), 
	.C0(n722), 
	.B0(n721), 
	.A1(n121), 
	.A0(n1575));
   OAI21XL U823 (.Y(n726), 
	.B0(n123), 
	.A1(n1592), 
	.A0(n32));
   NAND4X1 U824 (.Y(n1037), 
	.D(n1041), 
	.C(n1040), 
	.B(n1039), 
	.A(n1038));
   AOI21X1 U825 (.Y(n1040), 
	.B0(n179), 
	.A1(n1047), 
	.A0(n181));
   AOI211X1 U826 (.Y(n1041), 
	.C0(n1043), 
	.B0(n1042), 
	.A1(n118), 
	.A0(n190));
   OAI21XL U827 (.Y(n1047), 
	.B0(n120), 
	.A1(n207), 
	.A0(n33));
   NAND4X1 U828 (.Y(n454), 
	.D(n458), 
	.C(n457), 
	.B(n456), 
	.A(n455));
   AOI21X1 U829 (.Y(n457), 
	.B0(n1526), 
	.A1(n464), 
	.A0(n1528));
   AOI211X1 U830 (.Y(n458), 
	.C0(n460), 
	.B0(n459), 
	.A1(n115), 
	.A0(n1538));
   OAI21XL U831 (.Y(n464), 
	.B0(n117), 
	.A1(n1555), 
	.A0(n34));
   NAND4BXL U832 (.Y(n1349), 
	.D(n1353), 
	.C(n1352), 
	.B(n1284), 
	.AN(n1266));
   AOI221X1 U833 (.Y(n1353), 
	.C0(n1354), 
	.B1(n635), 
	.B0(n65), 
	.A1(n1102), 
	.A0(n50));
   AOI21XL U834 (.Y(n1354), 
	.B0(n23), 
	.A1(n1308), 
	.A0(n254));
   OAI21XL U835 (.Y(n1319), 
	.B0(n1320), 
	.A1(n247), 
	.A0(n262));
   OAI21XL U836 (.Y(n1320), 
	.B0(n1517), 
	.A1(n1502), 
	.A0(n635));
   OAI21XL U837 (.Y(n307), 
	.B0(n309), 
	.A1(sboxw[13]), 
	.A0(n308));
   AOI31X1 U838 (.Y(n309), 
	.B0(n276), 
	.A2(n49), 
	.A1(n1511), 
	.A0(n54));
   AOI211X1 U839 (.Y(n308), 
	.C0(n478), 
	.B0(n310), 
	.A1(n50), 
	.A0(n1509));
   INVX1 U840 (.Y(n478), 
	.A(n311));
   NAND4BXL U841 (.Y(n709), 
	.D(n712), 
	.C(n1587), 
	.B(n605), 
	.AN(n589));
   AOI211X1 U842 (.Y(n712), 
	.C0(n713), 
	.B0(n1562), 
	.A1(n30), 
	.A0(n1582));
   AOI21X1 U843 (.Y(n713), 
	.B0(n121), 
	.A1(n631), 
	.A0(n14));
   INVX1 U844 (.Y(n1562), 
	.A(n714));
   NAND4BXL U845 (.Y(n447), 
	.D(n450), 
	.C(n1548), 
	.B(n376), 
	.AN(n360));
   AOI211X1 U846 (.Y(n450), 
	.C0(n451), 
	.B0(n1558), 
	.A1(n31), 
	.A0(n1534));
   AOI21X1 U847 (.Y(n451), 
	.B0(n115), 
	.A1(n402), 
	.A0(n443));
   INVX1 U848 (.Y(n1558), 
	.A(n452));
   OAI211X1 U849 (.Y(n281), 
	.C0(n284), 
	.B0(n283), 
	.A1(n282), 
	.A0(n125));
   AOI31X1 U850 (.Y(n283), 
	.B0(n292), 
	.A2(n291), 
	.A1(n240), 
	.A0(n290));
   AOI222XL U851 (.Y(n284), 
	.C1(n247), 
	.C0(n273), 
	.B1(n25), 
	.B0(n286), 
	.A1(n285), 
	.A0(n153));
   NAND4X1 U852 (.Y(n285), 
	.D(n289), 
	.C(n288), 
	.B(n249), 
	.A(n287));
   AOI21XL U853 (.Y(n311), 
	.B0(n313), 
	.A1(n312), 
	.A0(n25));
   NAND4X1 U854 (.Y(n621), 
	.D(n633), 
	.C(n632), 
	.B(n631), 
	.A(n582));
   AOI22X1 U855 (.Y(n632), 
	.B1(n40), 
	.B0(n1575), 
	.A1(n4), 
	.A0(n634));
   AOI222X1 U856 (.Y(n633), 
	.C1(n576), 
	.C0(n1585), 
	.B1(n26), 
	.B0(n66), 
	.A1(n136), 
	.A0(n1593));
   NAND4X1 U857 (.Y(n975), 
	.D(n987), 
	.C(n986), 
	.B(n985), 
	.A(n936));
   AOI22X1 U858 (.Y(n986), 
	.B1(n38), 
	.B0(n190), 
	.A1(n15), 
	.A0(n988));
   AOI222X1 U859 (.Y(n987), 
	.C1(n930), 
	.C0(n195), 
	.B1(n27), 
	.B0(n203), 
	.A1(n148), 
	.A0(n56));
   NAND4X1 U860 (.Y(n392), 
	.D(n404), 
	.C(n403), 
	.B(n402), 
	.A(n353));
   AOI22X1 U861 (.Y(n403), 
	.B1(n39), 
	.B0(n1538), 
	.A1(n16), 
	.A0(n405));
   AOI222X1 U862 (.Y(n404), 
	.C1(n347), 
	.C0(n1543), 
	.B1(n28), 
	.B0(n1551), 
	.A1(n167), 
	.A0(n57));
   NAND4X1 U863 (.Y(n1169), 
	.D(n1180), 
	.C(n936), 
	.B(n1069), 
	.A(n1015));
   AOI32X1 U864 (.Y(n1180), 
	.B1(n33), 
	.B0(n1079), 
	.A2(n36), 
	.A1(n211), 
	.A0(n20));
   NAND4X1 U865 (.Y(n677), 
	.D(n688), 
	.C(n353), 
	.B(n486), 
	.A(n432));
   AOI32X1 U866 (.Y(n688), 
	.B1(n34), 
	.B0(n496), 
	.A2(n37), 
	.A1(n1559), 
	.A0(n21));
   NAND4X1 U867 (.Y(n867), 
	.D(n869), 
	.C(n868), 
	.B(n594), 
	.A(n717));
   AOI32X1 U868 (.Y(n868), 
	.B1(n123), 
	.B0(n772), 
	.A2(sboxw[24]), 
	.A1(n1594), 
	.A0(n1583));
   AOI222X1 U869 (.Y(n869), 
	.C1(n66), 
	.C0(n30), 
	.B1(n40), 
	.B0(n1576), 
	.A1(n26), 
	.A0(n63));
   NAND4X1 U870 (.Y(n1216), 
	.D(n1218), 
	.C(n1217), 
	.B(n948), 
	.A(n1038));
   AOI32X1 U871 (.Y(n1217), 
	.B1(n120), 
	.B0(n1093), 
	.A2(sboxw[16]), 
	.A1(n197), 
	.A0(n211));
   AOI222X1 U872 (.Y(n1218), 
	.C1(n203), 
	.C0(n29), 
	.B1(n38), 
	.B0(n202), 
	.A1(n27), 
	.A0(n64));
   NAND4X1 U873 (.Y(n1121), 
	.D(n1123), 
	.C(n1122), 
	.B(n365), 
	.A(n455));
   AOI32X1 U874 (.Y(n1122), 
	.B1(n117), 
	.B0(n510), 
	.A2(sboxw[0]), 
	.A1(n1545), 
	.A0(n1559));
   AOI222X1 U875 (.Y(n1123), 
	.C1(n1551), 
	.C0(n31), 
	.B1(n39), 
	.B0(n1550), 
	.A1(n28), 
	.A0(n1536));
   OAI21XL U876 (.Y(n896), 
	.B0(n898), 
	.A1(n129), 
	.A0(n897));
   AOI31X1 U877 (.Y(n898), 
	.B0(n1580), 
	.A2(n35), 
	.A1(n1592), 
	.A0(n1581));
   NOR4BX1 U878 (.Y(n897), 
	.D(n606), 
	.C(n1574), 
	.B(n900), 
	.AN(n899));
   AOI21X1 U879 (.Y(n899), 
	.B0(n627), 
	.A1(n1576), 
	.A0(n122));
   NAND4X1 U880 (.Y(n1446), 
	.D(n1459), 
	.C(n1289), 
	.B(n1384), 
	.A(n1334));
   AOI32X1 U881 (.Y(n1459), 
	.B1(n55), 
	.B0(n1509), 
	.A2(n124), 
	.A1(n1515), 
	.A0(n242));
   NAND4X1 U882 (.Y(n1369), 
	.D(n248), 
	.C(n298), 
	.B(n324), 
	.A(n1352));
   AOI21X1 U883 (.Y(n1140), 
	.B0(n143), 
	.A1(n952), 
	.A0(n18));
   AOI21X1 U884 (.Y(n529), 
	.B0(n159), 
	.A1(n369), 
	.A0(n19));
   NAND4X1 U885 (.Y(n255), 
	.D(n270), 
	.C(n269), 
	.B(n268), 
	.A(n267));
   AOI2BB2X1 U886 (.Y(n267), 
	.B1(n275), 
	.B0(n49), 
	.A1N(n277), 
	.A0N(n13));
   AOI31X1 U887 (.Y(n270), 
	.B0(n271), 
	.A2(n1502), 
	.A1(n1517), 
	.A0(sboxw[13]));
   AOI22XL U888 (.Y(n268), 
	.B1(n54), 
	.B0(n477), 
	.A1(n23), 
	.A0(n274));
   AOI21X1 U889 (.Y(n622), 
	.B0(n625), 
	.A1(n624), 
	.A0(n623));
   AOI222X1 U890 (.Y(n623), 
	.C1(n135), 
	.C0(n1576), 
	.B1(n11), 
	.B0(n629), 
	.A1(n136), 
	.A0(n1574));
   AOI211X1 U891 (.Y(n624), 
	.C0(n628), 
	.B0(n627), 
	.A1(n138), 
	.A0(n626));
   AOI21X1 U892 (.Y(n976), 
	.B0(n979), 
	.A1(n978), 
	.A0(n977));
   AOI222X1 U893 (.Y(n977), 
	.C1(sboxw[17]), 
	.C0(n202), 
	.B1(n8), 
	.B0(n983), 
	.A1(n146), 
	.A0(n198));
   AOI211X1 U894 (.Y(n978), 
	.C0(n982), 
	.B0(n981), 
	.A1(n151), 
	.A0(n980));
   AOI21X1 U895 (.Y(n393), 
	.B0(n396), 
	.A1(n395), 
	.A0(n394));
   AOI222X1 U896 (.Y(n394), 
	.C1(sboxw[1]), 
	.C0(n1550), 
	.B1(n7), 
	.B0(n400), 
	.A1(n167), 
	.A0(n1546));
   AOI211X1 U897 (.Y(n395), 
	.C0(n399), 
	.B0(n398), 
	.A1(n169), 
	.A0(n397));
   NAND4X1 U898 (.Y(n913), 
	.D(n939), 
	.C(n938), 
	.B(n937), 
	.A(n936));
   AOI221X1 U899 (.Y(n939), 
	.C0(n941), 
	.B1(n119), 
	.B0(n199), 
	.A1(n120), 
	.A0(n198));
   AOI21X1 U900 (.Y(n938), 
	.B0(n943), 
	.A1(n150), 
	.A0(n942));
   NAND4X1 U901 (.Y(n330), 
	.D(n356), 
	.C(n355), 
	.B(n354), 
	.A(n353));
   AOI221X1 U902 (.Y(n356), 
	.C0(n358), 
	.B1(n116), 
	.B0(n1547), 
	.A1(n117), 
	.A0(n1546));
   AOI21X1 U903 (.Y(n355), 
	.B0(n360), 
	.A1(n168), 
	.A0(n359));
   AOI21X1 U904 (.Y(n790), 
	.B0(n129), 
	.A1(n793), 
	.A0(n792));
   AOI222X1 U905 (.Y(n792), 
	.C1(n10), 
	.C0(n67), 
	.B1(n30), 
	.B0(n1586), 
	.A1(n1590), 
	.A0(n644));
   AOI211X1 U906 (.Y(n793), 
	.C0(n794), 
	.B0(n668), 
	.A1(n135), 
	.A0(n1575));
   AOI21X1 U907 (.Y(n794), 
	.B0(n26), 
	.A1(n631), 
	.A0(n643));
   AOI21X1 U908 (.Y(n1139), 
	.B0(n142), 
	.A1(n1142), 
	.A0(n1141));
   AOI222X1 U909 (.Y(n1141), 
	.C1(n6), 
	.C0(n199), 
	.B1(n29), 
	.B0(n61), 
	.A1(n204), 
	.A0(n998));
   AOI211X1 U910 (.Y(n1142), 
	.C0(n1143), 
	.B0(n1022), 
	.A1(sboxw[17]), 
	.A0(n190));
   AOI21X1 U911 (.Y(n1143), 
	.B0(n27), 
	.A1(n985), 
	.A0(n997));
   AOI21X1 U912 (.Y(n528), 
	.B0(n161), 
	.A1(n531), 
	.A0(n530));
   AOI222X1 U913 (.Y(n530), 
	.C1(n5), 
	.C0(n1547), 
	.B1(n31), 
	.B0(n62), 
	.A1(n1552), 
	.A0(n415));
   AOI211X1 U914 (.Y(n531), 
	.C0(n532), 
	.B0(n439), 
	.A1(sboxw[1]), 
	.A0(n1538));
   AOI21X1 U915 (.Y(n532), 
	.B0(n28), 
	.A1(n402), 
	.A0(n414));
   INVX1 U917 (.Y(n1061), 
	.A(n246));
   NAND3X1 U918 (.Y(n1184), 
	.C(n1187), 
	.B(n1186), 
	.A(n1185));
   NAND3X1 U919 (.Y(n1187), 
	.C(n181), 
	.B(n20), 
	.A(n8));
   NAND3X1 U920 (.Y(n692), 
	.C(n695), 
	.B(n694), 
	.A(n693));
   NAND3X1 U921 (.Y(n695), 
	.C(n1528), 
	.B(n21), 
	.A(n7));
   INVX1 U923 (.Y(n1506), 
	.A(n17));
   INVX1 U925 (.Y(n1586), 
	.A(n14));
   INVX1 U926 (.Y(n1536), 
	.A(n9));
   INVX1 U927 (.Y(n1507), 
	.A(n230));
   INVX1 U928 (.Y(n199), 
	.A(n18));
   INVX1 U929 (.Y(n1547), 
	.A(n19));
   INVX1 U930 (.Y(n1505), 
	.A(n1334));
   INVX1 U931 (.Y(n401), 
	.A(n1467));
   AOI221X1 U932 (.Y(n1467), 
	.C0(n1269), 
	.B1(n227), 
	.B0(n240), 
	.A1(n406), 
	.A0(n126));
   OAI2BB1X1 U933 (.Y(n1447), 
	.B0(n1453), 
	.A1N(n1452), 
	.A0N(n216));
   NAND4BXL U934 (.Y(n1452), 
	.D(n1457), 
	.C(n249), 
	.B(n1384), 
	.AN(n1456));
   OAI21XL U935 (.Y(n1453), 
	.B0(n219), 
	.A1(n1454), 
	.A0(n630));
   AOI21X1 U936 (.Y(n1457), 
	.B0(n1341), 
	.A1(n125), 
	.A0(n739));
   INVX1 U937 (.Y(n204), 
	.A(n20));
   INVX1 U938 (.Y(n1552), 
	.A(n21));
   INVX1 U939 (.Y(n203), 
	.A(n1));
   INVX1 U940 (.Y(n1551), 
	.A(n3));
   OAI222XL U944 (.Y(n607), 
	.C1(n129), 
	.C0(n612), 
	.B1(n611), 
	.B0(n130), 
	.A1(n597), 
	.A0(n599));
   AND3X2 U945 (.Y(n612), 
	.C(n615), 
	.B(n614), 
	.A(n613));
   AOI222X1 U946 (.Y(n613), 
	.C1(n1582), 
	.C0(n616), 
	.B1(n588), 
	.B0(n123), 
	.A1(n1574), 
	.A0(n32));
   INVX1 U947 (.Y(n175), 
	.A(n1156));
   AOI22X1 U948 (.Y(n1156), 
	.B1(n1158), 
	.B0(n176), 
	.A1(n1157), 
	.A0(n177));
   NAND4BXL U949 (.Y(n1157), 
	.D(n1162), 
	.C(n1069), 
	.B(n950), 
	.AN(n1161));
   NAND4X1 U950 (.Y(n1158), 
	.D(n1159), 
	.C(n1005), 
	.B(n999), 
	.A(n1089));
   INVX1 U951 (.Y(n137), 
	.A(n138));
   INVX1 U953 (.Y(n168), 
	.A(n169));
   INVX1 U958 (.Y(n163), 
	.A(n159));
   NAND2X1 U959 (.Y(n290), 
	.B(n242), 
	.A(n243));
   NOR2X1 U960 (.Y(n811), 
	.B(n772), 
	.A(n758));
   NOR2X1 U961 (.Y(n638), 
	.B(n604), 
	.A(n22));
   NOR2X1 U962 (.Y(n992), 
	.B(n958), 
	.A(n999));
   NOR2X1 U963 (.Y(n409), 
	.B(n375), 
	.A(n416));
   NOR2BX1 U964 (.Y(n789), 
	.B(n1592), 
	.AN(n577));
   NOR2BX1 U965 (.Y(n1138), 
	.B(n207), 
	.AN(n931));
   NOR2BX1 U966 (.Y(n527), 
	.B(n1555), 
	.AN(n348));
   NOR2X1 U967 (.Y(n606), 
	.B(n781), 
	.A(n11));
   NOR2X1 U968 (.Y(n983), 
	.B(n207), 
	.A(n211));
   NOR2X1 U969 (.Y(n400), 
	.B(n1555), 
	.A(n1559));
   NOR2X1 U970 (.Y(n1313), 
	.B(n1515), 
	.A(n1511));
   INVX1 U971 (.Y(n205), 
	.A(n1014));
   INVX1 U972 (.Y(n1553), 
	.A(n431));
   NOR2X1 U973 (.Y(n801), 
	.B(n2), 
	.A(n599));
   AOI211X1 U974 (.Y(n1390), 
	.C0(n58), 
	.B0(n275), 
	.A1(n1251), 
	.A0(n65));
   AOI211X1 U975 (.Y(n754), 
	.C0(n63), 
	.B0(n759), 
	.A1(n1594), 
	.A0(n30));
   AOI211X1 U976 (.Y(n1075), 
	.C0(n64), 
	.B0(n1080), 
	.A1(n197), 
	.A0(n29));
   AOI211X1 U977 (.Y(n492), 
	.C0(n1536), 
	.B0(n497), 
	.A1(n1545), 
	.A0(n31));
   OAI22X1 U978 (.Y(n759), 
	.B1(n2), 
	.B0(n135), 
	.A1(n136), 
	.A0(n1592));
   OAI22X1 U979 (.Y(n1080), 
	.B1(n20), 
	.B0(n147), 
	.A1(n148), 
	.A0(n207));
   OAI22X1 U980 (.Y(n497), 
	.B1(n21), 
	.B0(n166), 
	.A1(n167), 
	.A0(n1555));
   OAI22XL U981 (.Y(n1322), 
	.B1(n1333), 
	.B0(n247), 
	.A1(n254), 
	.A0(n54));
   NOR2XL U982 (.Y(n1335), 
	.B(n242), 
	.A(n318));
   NOR2XL U983 (.Y(n1270), 
	.B(n242), 
	.A(n1517));
   OAI211XL U984 (.Y(n1398), 
	.C0(n1400), 
	.B0(n1399), 
	.A1(n247), 
	.A0(n1374));
   AOI32X1 U985 (.Y(n1399), 
	.B1(n1495), 
	.B0(n124), 
	.A2(n645), 
	.A1(n1515), 
	.A0(n125));
   AOI21X1 U986 (.Y(n1400), 
	.B0(n1322), 
	.A1(n1061), 
	.A0(n65));
   OAI211X1 U987 (.Y(n1323), 
	.C0(n1338), 
	.B0(n1337), 
	.A1(n13), 
	.A0(n1336));
   AOI211X1 U988 (.Y(n1338), 
	.C0(n1341), 
	.B0(n1340), 
	.A1(n1339), 
	.A0(n291));
   AOI22X1 U989 (.Y(n1337), 
	.B1(n156), 
	.B0(n1344), 
	.A1(n1343), 
	.A0(n153));
   AOI2BB1X1 U990 (.Y(n1340), 
	.B0(n1342), 
	.A1N(n1270), 
	.A0N(n1513));
   OAI211X1 U991 (.Y(n890), 
	.C0(n595), 
	.B0(n605), 
	.A1(n642), 
	.A0(n891));
   NOR2X1 U992 (.Y(n232), 
	.B(n1516), 
	.A(n17));
   INVX1 U993 (.Y(n1596), 
	.A(n565));
   INVX1 U994 (.Y(n176), 
	.A(n919));
   INVX1 U995 (.Y(n1523), 
	.A(n336));
   NOR2X1 U996 (.Y(n778), 
	.B(n136), 
	.A(n781));
   NOR2X1 U997 (.Y(n1099), 
	.B(n148), 
	.A(n18));
   NOR2X1 U998 (.Y(n516), 
	.B(n167), 
	.A(n19));
   NAND2X1 U999 (.Y(n625), 
	.B(n1598), 
	.A(n129));
   NAND2X1 U1000 (.Y(n979), 
	.B(n174), 
	.A(n142));
   NAND2X1 U1001 (.Y(n396), 
	.B(n1521), 
	.A(n161));
   INVX1 U1002 (.Y(n219), 
	.A(n1330));
   AOI31X1 U1003 (.Y(n722), 
	.B0(n604), 
	.A2(n611), 
	.A1(n642), 
	.A0(n669));
   AOI31X1 U1004 (.Y(n815), 
	.B0(n725), 
	.A2(n811), 
	.A1(n1594), 
	.A0(n32));
   AOI21X1 U1005 (.Y(n237), 
	.B0(n1506), 
	.A1(n1507), 
	.A0(n1516));
   INVX1 U1006 (.Y(n1508), 
	.A(n1333));
   NOR2BX1 U1007 (.Y(n292), 
	.B(n1516), 
	.AN(n1335));
   INVX1 U1008 (.Y(n477), 
	.A(n1428));
   NOR2X1 U1009 (.Y(n841), 
	.B(sboxw[24]), 
	.A(n781));
   NOR2X1 U1010 (.Y(n662), 
	.B(n40), 
	.A(n634));
   NOR2X1 U1011 (.Y(n303), 
	.B(n1517), 
	.A(n1394));
   INVX1 U1012 (.Y(n1509), 
	.A(n1394));
   INVX1 U1013 (.Y(n1512), 
	.A(n314));
   OAI22X1 U1014 (.Y(n1408), 
	.B1(n314), 
	.B0(n50), 
	.A1(n1311), 
	.A0(n65));
   NOR2X1 U1015 (.Y(n581), 
	.B(n130), 
	.A(n14));
   INVX1 U1016 (.Y(n1513), 
	.A(n1361));
   NAND3X1 U1017 (.Y(n813), 
	.C(n811), 
	.B(n1594), 
	.A(n122));
   NAND3X1 U1018 (.Y(n1162), 
	.C(n1160), 
	.B(n197), 
	.A(n119));
   NAND3X1 U1019 (.Y(n551), 
	.C(n549), 
	.B(n1545), 
	.A(n116));
   NAND2X1 U1020 (.Y(n1352), 
	.B(n55), 
	.A(n239));
   NAND2X1 U1021 (.Y(n830), 
	.B(sboxw[24]), 
	.A(n758));
   NAND2X1 U1022 (.Y(n1179), 
	.B(n150), 
	.A(n1079));
   NAND2X1 U1023 (.Y(n687), 
	.B(sboxw[0]), 
	.A(n496));
   NAND2X1 U1024 (.Y(n566), 
	.B(n767), 
	.A(n14));
   AND2X2 U1025 (.Y(n50), 
	.B(n1517), 
	.A(n1516));
   NAND4X1 U1027 (.Y(n843), 
	.D(n847), 
	.C(n846), 
	.B(n643), 
	.A(n1587));
   AOI221X1 U1028 (.Y(n847), 
	.C0(n848), 
	.B1(n32), 
	.B0(n780), 
	.A1(n26), 
	.A0(n1574));
   AOI21X1 U1029 (.Y(n848), 
	.B0(n136), 
	.A1(n660), 
	.A0(n4));
   NAND2XL U1030 (.Y(n304), 
	.B(n23), 
	.A(n1335));
   AOI2BB2X1 U1031 (.Y(n872), 
	.B1(n759), 
	.B0(n1581), 
	.A1N(n587), 
	.A0N(n4));
   AOI2BB2X1 U1032 (.Y(n1221), 
	.B1(n1080), 
	.B0(n181), 
	.A1N(n941), 
	.A0N(n15));
   AOI2BB2X1 U1033 (.Y(n1126), 
	.B1(n497), 
	.B0(n1528), 
	.A1N(n358), 
	.A0N(n16));
   NAND2X1 U1034 (.Y(n714), 
	.B(n32), 
	.A(n588));
   AOI2BB2X1 U1035 (.Y(n874), 
	.B1(n876), 
	.B0(n130), 
	.A1N(n40), 
	.A0N(n600));
   OAI22X1 U1036 (.Y(n876), 
	.B1(n740), 
	.B0(n139), 
	.A1(n781), 
	.A0(n30));
   AOI2BB2X1 U1037 (.Y(n1223), 
	.B1(n1225), 
	.B0(sboxw[21]), 
	.A1N(n38), 
	.A0N(n954));
   OAI22XL U1038 (.Y(n1225), 
	.B1(n1), 
	.B0(n151), 
	.A1(n18), 
	.A0(n29));
   AOI2BB2X1 U1039 (.Y(n1128), 
	.B1(n1130), 
	.B0(n159), 
	.A1N(n39), 
	.A0N(n371));
   OAI22XL U1040 (.Y(n1130), 
	.B1(n3), 
	.B0(n169), 
	.A1(n19), 
	.A0(n31));
   OAI2BB2X1 U1041 (.Y(n777), 
	.B1(n767), 
	.B0(n30), 
	.A1N(n772), 
	.A0N(n122));
   OAI2BB2X1 U1042 (.Y(n1098), 
	.B1(n1088), 
	.B0(n29), 
	.A1N(n1093), 
	.A0N(n119));
   OAI2BB2X1 U1043 (.Y(n515), 
	.B1(n505), 
	.B0(n31), 
	.A1N(n510), 
	.A0N(n116));
   NAND2X1 U1044 (.Y(n836), 
	.B(n129), 
	.A(n626));
   NAND2X1 U1045 (.Y(n1297), 
	.B(n1516), 
	.A(n58));
   NAND4X1 U1046 (.Y(n820), 
	.D(n831), 
	.C(n582), 
	.B(n748), 
	.A(n661));
   AOI32X1 U1047 (.Y(n831), 
	.B1(n32), 
	.B0(n758), 
	.A2(n35), 
	.A1(n1583), 
	.A0(n2));
   AOI21X1 U1048 (.Y(n791), 
	.B0(sboxw[29]), 
	.A1(n598), 
	.A0(n781));
   NAND4X1 U1049 (.Y(n559), 
	.D(n585), 
	.C(n584), 
	.B(n583), 
	.A(n582));
   AOI221X1 U1050 (.Y(n585), 
	.C0(n587), 
	.B1(n122), 
	.B0(n67), 
	.A1(n123), 
	.A0(n1574));
   AOI21X1 U1051 (.Y(n584), 
	.B0(n589), 
	.A1(n137), 
	.A0(n588));
   NAND2X1 U1052 (.Y(n1435), 
	.B(n217), 
	.A(sboxw[13]));
   NAND2X1 U1053 (.Y(n1442), 
	.B(n217), 
	.A(n153));
   INVX1 U1054 (.Y(n1501), 
	.A(n298));
   OR2X2 U1055 (.Y(n1331), 
	.B(n50), 
	.A(n302));
   NAND3X1 U1056 (.Y(n835), 
	.C(n838), 
	.B(n837), 
	.A(n836));
   NAND3X1 U1057 (.Y(n838), 
	.C(n1581), 
	.B(n2), 
	.A(n11));
   NAND2X1 U1058 (.Y(n1427), 
	.B(n316), 
	.A(n17));
   INVX1 U1059 (.Y(n1590), 
	.A(n2));
   INVX1 U1060 (.Y(n1593), 
	.A(n22));
   OAI2BB1X1 U1063 (.Y(n1100), 
	.B0(n18), 
	.A1N(n1101), 
	.A0N(sboxw[16]));
   OAI2BB1X1 U1064 (.Y(n517), 
	.B0(n19), 
	.A1N(n518), 
	.A0N(n168));
   INVX1 U1065 (.Y(n519), 
	.A(n324));
   AND2X2 U1066 (.Y(n51), 
	.B(n2), 
	.A(n642));
   INVX1 U1067 (.Y(n730), 
	.A(n51));
   AND2X2 U1068 (.Y(n52), 
	.B(n20), 
	.A(n996));
   INVX1 U1069 (.Y(n1051), 
	.A(n52));
   AND2X2 U1070 (.Y(n53), 
	.B(n21), 
	.A(n9));
   INVX1 U1071 (.Y(n468), 
	.A(n53));
   INVX1 U1072 (.Y(n672), 
	.A(n1328));
   OAI21XL U1073 (.Y(n1328), 
	.B0(n237), 
	.A1(n1321), 
	.A0(n243));
   NOR2X1 U1074 (.Y(n629), 
	.B(n1592), 
	.A(n1583));
   INVX1 U1075 (.Y(n1588), 
	.A(n660));
   INVX1 U1076 (.Y(n1597), 
	.A(n657));
   INVX1 U1077 (.Y(n177), 
	.A(n1011));
   INVX1 U1078 (.Y(n1524), 
	.A(n428));
   NAND2X1 U1079 (.Y(n262), 
	.B(n1251), 
	.A(n1515));
   INVX1 U1080 (.Y(n218), 
	.A(n223));
   OAI22XL U1081 (.Y(n1409), 
	.B1(n1333), 
	.B0(n25), 
	.A1(n247), 
	.A0(n230));
   NAND2X1 U1082 (.Y(n1401), 
	.B(n65), 
	.A(n312));
   AOI2BB2XL U1083 (.Y(n260), 
	.B1(n24), 
	.B0(n1512), 
	.A1N(n1517), 
	.A0N(n262));
   INVX1 U1084 (.Y(n214), 
	.A(n1346));
   OAI2BB1X1 U1085 (.Y(n779), 
	.B0(n781), 
	.A1N(n780), 
	.A0N(sboxw[24]));
   INVX1 U1086 (.Y(n1599), 
	.A(n555));
   INVX1 U1087 (.Y(n172), 
	.A(n909));
   INVX1 U1088 (.Y(n1519), 
	.A(n326));
   INVX1 U1089 (.Y(n213), 
	.A(n1258));
   OAI222XL U1090 (.Y(new_sboxw[18]), 
	.C1(n1167), 
	.C0(sboxw[23]), 
	.B1(n911), 
	.B0(n1166), 
	.A1(n909), 
	.A0(n1165));
   AOI221X1 U1091 (.Y(n1165), 
	.C0(n1193), 
	.B1(n142), 
	.B0(n1192), 
	.A1(n1191), 
	.A0(n143));
   AOI221X1 U1092 (.Y(n1166), 
	.C0(n1184), 
	.B1(n1183), 
	.B0(sboxw[21]), 
	.A1(n148), 
	.A0(n1138));
   AOI221X1 U1093 (.Y(n1167), 
	.C0(n1170), 
	.B1(n1169), 
	.B0(n176), 
	.A1(n1168), 
	.A0(n974));
   OAI222XL U1094 (.Y(new_sboxw[23]), 
	.C1(n912), 
	.C0(sboxw[23]), 
	.B1(n911), 
	.B0(n910), 
	.A1(n909), 
	.A0(n908));
   NOR4X1 U1095 (.Y(n910), 
	.D(n947), 
	.C(n946), 
	.B(n945), 
	.A(n944));
   AOI211X1 U1096 (.Y(n908), 
	.C0(n962), 
	.B0(n961), 
	.A1(n199), 
	.A0(n933));
   AOI211X1 U1097 (.Y(n912), 
	.C0(n915), 
	.B0(n914), 
	.A1(n913), 
	.A0(n177));
   OAI222XL U1098 (.Y(new_sboxw[21]), 
	.C1(n909), 
	.C0(n1029), 
	.B1(n1028), 
	.B0(sboxw[23]), 
	.A1(n911), 
	.A0(n1027));
   AOI222X1 U1099 (.Y(n1029), 
	.C1(n1032), 
	.C0(n181), 
	.B1(n142), 
	.B0(n1031), 
	.A1(n1030), 
	.A0(sboxw[21]));
   NOR4BBX1 U1100 (.Y(n1027), 
	.D(n921), 
	.C(n932), 
	.BN(n1057), 
	.AN(n1056));
   AOI22X1 U1101 (.Y(n1028), 
	.B1(n174), 
	.B0(n1037), 
	.A1(n1036), 
	.A0(sboxw[22]));
   OAI222XL U1102 (.Y(new_sboxw[2]), 
	.C1(n675), 
	.C0(sboxw[7]), 
	.B1(n328), 
	.B0(n674), 
	.A1(n326), 
	.A0(n673));
   AOI221X1 U1103 (.Y(n673), 
	.C0(n701), 
	.B1(n160), 
	.B0(n700), 
	.A1(n699), 
	.A0(sboxw[5]));
   AOI221X1 U1104 (.Y(n674), 
	.C0(n692), 
	.B1(n691), 
	.B0(sboxw[5]), 
	.A1(n167), 
	.A0(n527));
   AOI221X1 U1105 (.Y(n675), 
	.C0(n678), 
	.B1(n677), 
	.B0(n1523), 
	.A1(n676), 
	.A0(n391));
   OAI222XL U1106 (.Y(new_sboxw[7]), 
	.C1(n329), 
	.C0(sboxw[7]), 
	.B1(n328), 
	.B0(n327), 
	.A1(n326), 
	.A0(n325));
   NOR4X1 U1107 (.Y(n327), 
	.D(n364), 
	.C(n363), 
	.B(n362), 
	.A(n361));
   AOI211X1 U1108 (.Y(n325), 
	.C0(n379), 
	.B0(n378), 
	.A1(n1547), 
	.A0(n350));
   AOI211X1 U1109 (.Y(n329), 
	.C0(n332), 
	.B0(n331), 
	.A1(n330), 
	.A0(n1524));
   OAI222X1 U1110 (.Y(new_sboxw[5]), 
	.C1(n326), 
	.C0(n446), 
	.B1(n445), 
	.B0(sboxw[7]), 
	.A1(n328), 
	.A0(n444));
   AOI222X1 U1111 (.Y(n446), 
	.C1(n449), 
	.C0(n1528), 
	.B1(n160), 
	.B0(n448), 
	.A1(n447), 
	.A0(sboxw[5]));
   NOR4BBX1 U1112 (.Y(n444), 
	.D(n338), 
	.C(n349), 
	.BN(n474), 
	.AN(n473));
   AOI22X1 U1113 (.Y(n445), 
	.B1(n1521), 
	.B0(n454), 
	.A1(n453), 
	.A0(sboxw[6]));
   OAI222XL U1114 (.Y(new_sboxw[26]), 
	.C1(n818), 
	.C0(sboxw[31]), 
	.B1(n557), 
	.B0(n817), 
	.A1(n555), 
	.A0(n816));
   AOI221X1 U1115 (.Y(n816), 
	.C0(n844), 
	.B1(n128), 
	.B0(n843), 
	.A1(n842), 
	.A0(n130));
   AOI221X1 U1116 (.Y(n817), 
	.C0(n835), 
	.B1(n834), 
	.B0(n130), 
	.A1(n136), 
	.A0(n789));
   AOI221X1 U1117 (.Y(n818), 
	.C0(n821), 
	.B1(n820), 
	.B0(n1596), 
	.A1(n819), 
	.A0(n620));
   OAI22X1 U1118 (.Y(new_sboxw[16]), 
	.B1(n1227), 
	.B0(sboxw[23]), 
	.A1(n171), 
	.A0(n1226));
   AOI222X1 U1119 (.Y(n1226), 
	.C1(n1245), 
	.C0(sboxw[22]), 
	.B1(n1244), 
	.B0(n176), 
	.A1(n174), 
	.A0(n1243));
   AOI22X1 U1120 (.Y(n1227), 
	.B1(n174), 
	.B0(n1229), 
	.A1(n1228), 
	.A0(sboxw[22]));
   OAI221XL U1121 (.Y(n1244), 
	.C0(n952), 
	.B1(n996), 
	.B0(n1240), 
	.A1(n970), 
	.A0(n1));
   OAI22X1 U1122 (.Y(new_sboxw[0]), 
	.B1(n1471), 
	.B0(sboxw[7]), 
	.A1(n1518), 
	.A0(n1470));
   AOI222X1 U1123 (.Y(n1470), 
	.C1(n1489), 
	.C0(sboxw[6]), 
	.B1(n1488), 
	.B0(n1523), 
	.A1(n1521), 
	.A0(n1487));
   AOI22X1 U1124 (.Y(n1471), 
	.B1(n1521), 
	.B0(n1473), 
	.A1(n1472), 
	.A0(sboxw[6]));
   OAI221XL U1125 (.Y(n1488), 
	.C0(n369), 
	.B1(n9), 
	.B0(n1484), 
	.A1(n387), 
	.A0(n3));
   NAND2X1 U1126 (.Y(n643), 
	.B(sboxw[26]), 
	.A(n1591));
   NAND2X1 U1127 (.Y(n997), 
	.B(sboxw[18]), 
	.A(n196));
   NAND2X1 U1128 (.Y(n414), 
	.B(sboxw[2]), 
	.A(n1544));
   OAI2BB2X1 U1129 (.Y(new_sboxw[17]), 
	.B1(n1198), 
	.B0(sboxw[23]), 
	.A1N(n1199), 
	.A0N(sboxw[23]));
   AOI222X1 U1130 (.Y(n1198), 
	.C1(n1216), 
	.C0(n176), 
	.B1(n1215), 
	.B0(n177), 
	.A1(n174), 
	.A0(n1214));
   OAI221XL U1131 (.Y(n1199), 
	.C0(n1202), 
	.B1(n1201), 
	.B0(sboxw[22]), 
	.A1(n919), 
	.A0(n1200));
   NAND4X1 U1132 (.Y(n1214), 
	.D(n1224), 
	.C(n1223), 
	.B(n1222), 
	.A(n1221));
   OAI2BB2X1 U1133 (.Y(new_sboxw[1]), 
	.B1(n1103), 
	.B0(sboxw[7]), 
	.A1N(n1104), 
	.A0N(sboxw[7]));
   AOI222X1 U1134 (.Y(n1103), 
	.C1(n1121), 
	.C0(n1523), 
	.B1(n1120), 
	.B0(n1524), 
	.A1(n1521), 
	.A0(n1119));
   OAI221XL U1135 (.Y(n1104), 
	.C0(n1107), 
	.B1(n1106), 
	.B0(sboxw[6]), 
	.A1(n336), 
	.A0(n1105));
   NAND4X1 U1136 (.Y(n1119), 
	.D(n1129), 
	.C(n1128), 
	.B(n1127), 
	.A(n1126));
   INVX1 U1137 (.Y(n1594), 
	.A(sboxw[28]));
   INVX1 U1138 (.Y(n1545), 
	.A(sboxw[4]));
   INVX1 U1139 (.Y(n197), 
	.A(sboxw[20]));
   OAI21XL U1140 (.Y(new_sboxw[20]), 
	.B0(n1065), 
	.A1(n171), 
	.A0(n1064));
   OAI2BB1X1 U1141 (.Y(n1065), 
	.B0(n171), 
	.A1N(n1067), 
	.A0N(n1066));
   AOI222X1 U1142 (.Y(n1064), 
	.C1(n1085), 
	.C0(n974), 
	.B1(n1084), 
	.B0(n173), 
	.A1(n1083), 
	.A0(sboxw[22]));
   AOI22X1 U1143 (.Y(n1067), 
	.B1(n1068), 
	.B0(n173), 
	.A1(n992), 
	.A0(n33));
   OAI21XL U1144 (.Y(new_sboxw[4]), 
	.B0(n482), 
	.A1(n1518), 
	.A0(n481));
   OAI2BB1X1 U1145 (.Y(n482), 
	.B0(n1518), 
	.A1N(n484), 
	.A0N(n483));
   AOI222X1 U1146 (.Y(n481), 
	.C1(n502), 
	.C0(n391), 
	.B1(n501), 
	.B0(n1520), 
	.A1(n500), 
	.A0(sboxw[6]));
   AOI22X1 U1147 (.Y(n484), 
	.B1(n485), 
	.B0(n1520), 
	.A1(n409), 
	.A0(n34));
   OAI21XL U1148 (.Y(new_sboxw[19]), 
	.B0(n1132), 
	.A1(n1131), 
	.A0(sboxw[23]));
   AOI211X1 U1149 (.Y(n1131), 
	.C0(n1152), 
	.B0(n175), 
	.A1(n1151), 
	.A0(n974));
   AOI21X1 U1150 (.Y(n1132), 
	.B0(n1134), 
	.A1(n1133), 
	.A0(n172));
   OAI221XL U1151 (.Y(n1151), 
	.C0(n1164), 
	.B1(n6), 
	.B0(n18), 
	.A1(n997), 
	.A0(n151));
   OAI21XL U1152 (.Y(new_sboxw[3]), 
	.B0(n521), 
	.A1(n520), 
	.A0(sboxw[7]));
   AOI211X1 U1153 (.Y(n520), 
	.C0(n541), 
	.B0(n1522), 
	.A1(n540), 
	.A0(n391));
   AOI21X1 U1154 (.Y(n521), 
	.B0(n523), 
	.A1(n522), 
	.A0(n1519));
   OAI221XL U1155 (.Y(n540), 
	.C0(n553), 
	.B1(n5), 
	.B0(n19), 
	.A1(n414), 
	.A0(n170));
   OAI22X1 U1156 (.Y(new_sboxw[24]), 
	.B1(n878), 
	.B0(sboxw[31]), 
	.A1(n1600), 
	.A0(n877));
   AOI222X1 U1157 (.Y(n877), 
	.C1(n896), 
	.C0(sboxw[30]), 
	.B1(n895), 
	.B0(n1596), 
	.A1(n1598), 
	.A0(n894));
   AOI22X1 U1158 (.Y(n878), 
	.B1(n1598), 
	.B0(n880), 
	.A1(n879), 
	.A0(sboxw[30]));
   OAI221XL U1159 (.Y(n895), 
	.C0(n598), 
	.B1(n642), 
	.B0(n891), 
	.A1(n616), 
	.A0(n740));
   OAI2BB2X1 U1160 (.Y(new_sboxw[25]), 
	.B1(n849), 
	.B0(sboxw[31]), 
	.A1N(n850), 
	.A0N(sboxw[31]));
   AOI222X1 U1161 (.Y(n849), 
	.C1(n867), 
	.C0(n1596), 
	.B1(n866), 
	.B0(n1597), 
	.A1(n1598), 
	.A0(n865));
   OAI221XL U1162 (.Y(n850), 
	.C0(n853), 
	.B1(n852), 
	.B0(sboxw[30]), 
	.A1(n565), 
	.A0(n851));
   NAND4X1 U1163 (.Y(n865), 
	.D(n875), 
	.C(n874), 
	.B(n873), 
	.A(n872));
   AOI32X1 U1164 (.Y(n853), 
	.B1(n854), 
	.B0(n1597), 
	.A2(n1577), 
	.A1(n123), 
	.A0(sboxw[30]));
   OAI221XL U1165 (.Y(n854), 
	.C0(n855), 
	.B1(n123), 
	.B0(n22), 
	.A1(n740), 
	.A0(n30));
   AOI211X1 U1166 (.Y(n855), 
	.C0(n1566), 
	.B0(n778), 
	.A1(n576), 
	.A0(n1586));
   INVX1 U1167 (.Y(n1566), 
	.A(n733));
   AOI32X1 U1168 (.Y(n1202), 
	.B1(n1203), 
	.B0(n177), 
	.A2(n184), 
	.A1(n120), 
	.A0(sboxw[22]));
   OAI221XL U1169 (.Y(n1203), 
	.C0(n1204), 
	.B1(n120), 
	.B0(n999), 
	.A1(n1), 
	.A0(n29));
   AOI211X1 U1170 (.Y(n1204), 
	.C0(n191), 
	.B0(n1099), 
	.A1(n930), 
	.A0(n61));
   INVX1 U1171 (.Y(n191), 
	.A(n1054));
   AOI32X1 U1172 (.Y(n1107), 
	.B1(n1108), 
	.B0(n1524), 
	.A2(n1531), 
	.A1(n117), 
	.A0(sboxw[6]));
   OAI221XL U1173 (.Y(n1108), 
	.C0(n1109), 
	.B1(n117), 
	.B0(n416), 
	.A1(n3), 
	.A0(n31));
   AOI211X1 U1174 (.Y(n1109), 
	.C0(n1539), 
	.B0(n516), 
	.A1(n347), 
	.A0(n62));
   INVX1 U1175 (.Y(n1539), 
	.A(n471));
   AOI31X1 U1176 (.Y(n914), 
	.B0(sboxw[22]), 
	.A2(n924), 
	.A1(n923), 
	.A0(n922));
   AOI2BB2X1 U1177 (.Y(n922), 
	.B1(n56), 
	.B0(n933), 
	.A1N(n29), 
	.A0N(n934));
   AOI31X1 U1178 (.Y(n923), 
	.B0(n932), 
	.A2(n931), 
	.A1(n207), 
	.A0(n930));
   AOI221X1 U1179 (.Y(n924), 
	.C0(n926), 
	.B1(n119), 
	.B0(n184), 
	.A1(sboxw[17]), 
	.A0(n198));
   AOI31X1 U1180 (.Y(n331), 
	.B0(sboxw[6]), 
	.A2(n341), 
	.A1(n340), 
	.A0(n339));
   AOI2BB2X1 U1181 (.Y(n339), 
	.B1(n57), 
	.B0(n350), 
	.A1N(n31), 
	.A0N(n351));
   AOI31X1 U1182 (.Y(n340), 
	.B0(n349), 
	.A2(n348), 
	.A1(n1555), 
	.A0(n347));
   AOI221X1 U1183 (.Y(n341), 
	.C0(n343), 
	.B1(n116), 
	.B0(n1531), 
	.A1(sboxw[1]), 
	.A0(n1546));
   AOI22X1 U1184 (.Y(n1066), 
	.B1(n1073), 
	.B0(sboxw[22]), 
	.A1(n1072), 
	.A0(n974));
   OAI221XL U1185 (.Y(n1072), 
	.C0(n1082), 
	.B1(n15), 
	.B0(n29), 
	.A1(n996), 
	.A0(n27));
   OAI222XL U1186 (.Y(n1073), 
	.C1(n142), 
	.C0(n1076), 
	.B1(n953), 
	.B0(n1075), 
	.A1(n1074), 
	.A0(sboxw[21]));
   AOI211X1 U1187 (.Y(n1082), 
	.C0(n943), 
	.B0(n61), 
	.A1(sboxw[17]), 
	.A0(n983));
   OAI21XL U1188 (.Y(new_sboxw[27]), 
	.B0(n783), 
	.A1(n782), 
	.A0(sboxw[31]));
   AOI211X1 U1189 (.Y(n782), 
	.C0(n803), 
	.B0(n1564), 
	.A1(n802), 
	.A0(n620));
   AOI21X1 U1190 (.Y(n783), 
	.B0(n785), 
	.A1(n784), 
	.A0(n1599));
   OAI221XL U1191 (.Y(n802), 
	.C0(n815), 
	.B1(n10), 
	.B0(n781), 
	.A1(n643), 
	.A0(n138));
   OAI222X1 U1192 (.Y(new_sboxw[13]), 
	.C1(n1258), 
	.C0(n1348), 
	.B1(n1347), 
	.B0(sboxw[15]), 
	.A1(n1346), 
	.A0(n1345));
   AOI222X1 U1193 (.Y(n1348), 
	.C1(n1351), 
	.C0(n49), 
	.B1(n156), 
	.B0(n1350), 
	.A1(n1349), 
	.A0(n153));
   NOR4BX1 U1194 (.Y(n1345), 
	.D(n1286), 
	.C(n263), 
	.B(n1373), 
	.AN(n1372));
   AOI22X1 U1195 (.Y(n1347), 
	.B1(n217), 
	.B0(n1356), 
	.A1(n1355), 
	.A0(sboxw[14]));
   OAI222XL U1196 (.Y(new_sboxw[10]), 
	.C1(n1445), 
	.C0(sboxw[15]), 
	.B1(n1346), 
	.B0(n1444), 
	.A1(n1258), 
	.A0(n1443));
   NOR4X1 U1197 (.Y(n1444), 
	.D(n286), 
	.C(n292), 
	.B(n1461), 
	.A(n1460));
   AOI221X1 U1198 (.Y(n1443), 
	.C0(n401), 
	.B1(n156), 
	.B0(n1466), 
	.A1(n1465), 
	.A0(n153));
   AOI211X1 U1199 (.Y(n1445), 
	.C0(n1448), 
	.B0(n1447), 
	.A1(n1446), 
	.A0(n218));
   OAI221XL U1200 (.Y(new_sboxw[15]), 
	.C0(n1260), 
	.B1(n1259), 
	.B0(sboxw[15]), 
	.A1(n1258), 
	.A0(n1257));
   OAI21XL U1201 (.Y(n1260), 
	.B0(n214), 
	.A1(n1262), 
	.A0(n1261));
   AOI211X1 U1202 (.Y(n1259), 
	.C0(n1273), 
	.B0(n1272), 
	.A1(n1271), 
	.A0(n219));
   AOI211X1 U1203 (.Y(n1257), 
	.C0(n1294), 
	.B0(n1293), 
	.A1(n1506), 
	.A0(n1287));
   OAI222XL U1204 (.Y(new_sboxw[29]), 
	.C1(n555), 
	.C0(n708), 
	.B1(n707), 
	.B0(sboxw[31]), 
	.A1(n557), 
	.A0(n706));
   AOI222X1 U1205 (.Y(n708), 
	.C1(n711), 
	.C0(n1581), 
	.B1(n128), 
	.B0(n710), 
	.A1(n709), 
	.A0(n130));
   NOR4BBX1 U1206 (.Y(n706), 
	.D(n567), 
	.C(n578), 
	.BN(n736), 
	.AN(n735));
   AOI22X1 U1207 (.Y(n707), 
	.B1(n1598), 
	.B0(n716), 
	.A1(n715), 
	.A0(sboxw[30]));
   OAI222XL U1208 (.Y(new_sboxw[31]), 
	.C1(n558), 
	.C0(sboxw[31]), 
	.B1(n557), 
	.B0(n556), 
	.A1(n555), 
	.A0(n554));
   NOR4X1 U1209 (.Y(n556), 
	.D(n593), 
	.C(n592), 
	.B(n591), 
	.A(n590));
   AOI211X1 U1210 (.Y(n554), 
	.C0(n608), 
	.B0(n607), 
	.A1(n67), 
	.A0(n579));
   AOI211X1 U1211 (.Y(n558), 
	.C0(n561), 
	.B0(n560), 
	.A1(n559), 
	.A0(n1597));
   OAI22X1 U1212 (.Y(new_sboxw[22]), 
	.B1(n171), 
	.B0(n972), 
	.A1(n971), 
	.A0(sboxw[23]));
   AOI211X1 U1213 (.Y(n971), 
	.C0(n1004), 
	.B0(n1003), 
	.A1(n174), 
	.A0(n1002));
   AOI221X1 U1214 (.Y(n972), 
	.C0(n976), 
	.B1(n975), 
	.B0(n974), 
	.A1(n973), 
	.A0(sboxw[22]));
   OAI211X1 U1215 (.Y(n1002), 
	.C0(n1019), 
	.B0(n1018), 
	.A1(n15), 
	.A0(n1017));
   OAI22X1 U1216 (.Y(new_sboxw[6]), 
	.B1(n1518), 
	.B0(n389), 
	.A1(n388), 
	.A0(sboxw[7]));
   AOI211X1 U1217 (.Y(n388), 
	.C0(n421), 
	.B0(n420), 
	.A1(n1521), 
	.A0(n419));
   AOI221X1 U1218 (.Y(n389), 
	.C0(n393), 
	.B1(n392), 
	.B0(n391), 
	.A1(n390), 
	.A0(sboxw[6]));
   OAI211X1 U1219 (.Y(n419), 
	.C0(n436), 
	.B0(n435), 
	.A1(n16), 
	.A0(n434));
   OAI22X1 U1220 (.Y(new_sboxw[14]), 
	.B1(n212), 
	.B0(n1304), 
	.A1(n1303), 
	.A0(sboxw[15]));
   AOI211X1 U1221 (.Y(n1303), 
	.C0(n1325), 
	.B0(n1324), 
	.A1(n217), 
	.A0(n1323));
   AOI222X1 U1222 (.Y(n1304), 
	.C1(n1307), 
	.C0(n215), 
	.B1(n1306), 
	.B0(n216), 
	.A1(n1305), 
	.A0(sboxw[14]));
   AOI31X1 U1223 (.Y(n1325), 
	.B0(n223), 
	.A2(n672), 
	.A1(n1327), 
	.A0(n1326));
   OAI22X1 U1224 (.Y(new_sboxw[8]), 
	.B1(n279), 
	.B0(sboxw[15]), 
	.A1(n212), 
	.A0(n278));
   AOI22X1 U1225 (.Y(n279), 
	.B1(n217), 
	.B0(n281), 
	.A1(n280), 
	.A0(sboxw[14]));
   AOI222X1 U1226 (.Y(n278), 
	.C1(n307), 
	.C0(sboxw[14]), 
	.B1(n306), 
	.B0(n218), 
	.A1(n217), 
	.A0(n305));
   OAI211X1 U1227 (.Y(n280), 
	.C0(n294), 
	.B0(n293), 
	.A1(n282), 
	.A0(n1517));
   OAI2BB2X1 U1228 (.Y(new_sboxw[9]), 
	.B1(n220), 
	.B0(sboxw[15]), 
	.A1N(n221), 
	.A0N(sboxw[15]));
   AOI222X1 U1229 (.Y(n220), 
	.C1(n257), 
	.C0(n218), 
	.B1(n256), 
	.B0(n219), 
	.A1(n217), 
	.A0(n255));
   OAI221XL U1230 (.Y(n221), 
	.C0(n225), 
	.B1(n224), 
	.B0(sboxw[14]), 
	.A1(n223), 
	.A0(n222));
   NAND4X1 U1231 (.Y(n257), 
	.D(n261), 
	.C(n260), 
	.B(n259), 
	.A(n258));
   INVX1 U1232 (.Y(n1251), 
	.A(sboxw[12]));
   OAI21X1 U1233 (.Y(new_sboxw[12]), 
	.B0(n1380), 
	.A1(n212), 
	.A0(n1379));
   OAI2BB1X1 U1234 (.Y(n1380), 
	.B0(n212), 
	.A1N(n1382), 
	.A0N(n1381));
   AOI222X1 U1235 (.Y(n1379), 
	.C1(n1398), 
	.C0(n215), 
	.B1(n1397), 
	.B0(n216), 
	.A1(n1396), 
	.A0(sboxw[14]));
   AOI22X1 U1236 (.Y(n1382), 
	.B1(n1383), 
	.B0(n216), 
	.A1(n274), 
	.A0(n55));
   OAI21XL U1237 (.Y(new_sboxw[11]), 
	.B0(n1411), 
	.A1(n1410), 
	.A0(sboxw[15]));
   AOI211X1 U1238 (.Y(n1410), 
	.C0(n1431), 
	.B0(n1430), 
	.A1(n1429), 
	.A0(n215));
   AOI22X1 U1239 (.Y(n1411), 
	.B1(n1413), 
	.B0(n213), 
	.A1(n1412), 
	.A0(n214));
   OAI221XL U1240 (.Y(n1429), 
	.C0(n1441), 
	.B1(n17), 
	.B0(n25), 
	.A1(n1517), 
	.A0(n246));
   NAND2X1 U1241 (.Y(n230), 
	.B(sboxw[11]), 
	.A(sboxw[12]));
   NAND2X1 U1242 (.Y(n246), 
	.B(n1102), 
	.A(sboxw[10]));
   NOR2X1 U1243 (.Y(n1079), 
	.B(sboxw[19]), 
	.A(n211));
   NOR2X1 U1244 (.Y(n496), 
	.B(sboxw[3]), 
	.A(n1559));
   AOI222X1 U1245 (.Y(n300), 
	.C1(n1503), 
	.C0(n65), 
	.B1(n124), 
	.B0(n301), 
	.A1(n1102), 
	.A0(sboxw[8]));
   NAND4X1 U1246 (.Y(n1084), 
	.D(n1092), 
	.C(n1091), 
	.B(n1090), 
	.A(n1089));
   NAND3X1 U1247 (.Y(n1091), 
	.C(n52), 
	.B(n118), 
	.A(sboxw[18]));
   AOI222X1 U1248 (.Y(n1092), 
	.C1(n36), 
	.C0(n190), 
	.B1(sboxw[17]), 
	.B0(n1093), 
	.A1(n119), 
	.A0(n61));
   AOI22X1 U1249 (.Y(n746), 
	.B1(n747), 
	.B0(n1595), 
	.A1(n638), 
	.A0(n32));
   NAND4X1 U1250 (.Y(n747), 
	.D(n750), 
	.C(n749), 
	.B(n1587), 
	.A(n748));
   NAND3X1 U1251 (.Y(n749), 
	.C(sboxw[26]), 
	.B(n121), 
	.A(n730));
   AOI222X1 U1252 (.Y(n750), 
	.C1(n32), 
	.C0(n1574), 
	.B1(n40), 
	.B0(n626), 
	.A1(n10), 
	.A0(n1575));
   NAND4X1 U1253 (.Y(n1068), 
	.D(n1071), 
	.C(n1070), 
	.B(n200), 
	.A(n1069));
   NAND3X1 U1254 (.Y(n1070), 
	.C(sboxw[18]), 
	.B(n118), 
	.A(n1051));
   AOI222X1 U1255 (.Y(n1071), 
	.C1(n33), 
	.C0(n198), 
	.B1(n38), 
	.B0(n980), 
	.A1(n6), 
	.A0(n190));
   NAND4X1 U1256 (.Y(n485), 
	.D(n488), 
	.C(n487), 
	.B(n1548), 
	.A(n486));
   NAND3X1 U1257 (.Y(n487), 
	.C(sboxw[2]), 
	.B(n115), 
	.A(n468));
   AOI222X1 U1258 (.Y(n488), 
	.C1(n34), 
	.C0(n1546), 
	.B1(n39), 
	.B0(n397), 
	.A1(n5), 
	.A0(n1538));
   OAI222XL U1259 (.Y(n1454), 
	.C1(n24), 
	.C0(n242), 
	.B1(n1308), 
	.B0(sboxw[9]), 
	.A1(n254), 
	.A0(n127));
   AOI22X1 U1260 (.Y(n644), 
	.B1(n32), 
	.B0(sboxw[26]), 
	.A1(n139), 
	.A0(n1583));
   AOI22X1 U1261 (.Y(n998), 
	.B1(n33), 
	.B0(sboxw[18]), 
	.A1(n151), 
	.A0(n211));
   AOI22X1 U1262 (.Y(n415), 
	.B1(n34), 
	.B0(sboxw[2]), 
	.A1(n169), 
	.A0(n1559));
   OAI222XL U1263 (.Y(n1396), 
	.C1(n1406), 
	.C0(n153), 
	.B1(n1342), 
	.B0(n1405), 
	.A1(sboxw[13]), 
	.A0(n1404));
   AOI21X1 U1264 (.Y(n1405), 
	.B0(n571), 
	.A1(n25), 
	.A0(n1102));
   AOI211X1 U1265 (.Y(n1404), 
	.C0(n1506), 
	.B0(n1409), 
	.A1(sboxw[8]), 
	.A0(n301));
   AOI211X1 U1266 (.Y(n1406), 
	.C0(n1408), 
	.B0(n1407), 
	.A1(n1516), 
	.A0(n739));
   AOI31X1 U1267 (.Y(n1448), 
	.B0(n1442), 
	.A2(n1451), 
	.A1(n1450), 
	.A0(n1449));
   AOI21X1 U1268 (.Y(n1450), 
	.B0(n1505), 
	.A1(n50), 
	.A0(n312));
   AOI22X1 U1269 (.Y(n1449), 
	.B1(sboxw[10]), 
	.B0(n1513), 
	.A1(n125), 
	.A0(n1509));
   AOI222XL U1270 (.Y(n1451), 
	.C1(n24), 
	.C0(n635), 
	.B1(n1516), 
	.B0(n1495), 
	.A1(n23), 
	.A0(n1102));
   AOI222X1 U1271 (.Y(n860), 
	.C1(n136), 
	.C0(n1588), 
	.B1(n35), 
	.B0(n588), 
	.A1(sboxw[26]), 
	.A0(n1568));
   AOI222X1 U1272 (.Y(n1209), 
	.C1(n148), 
	.C0(n205), 
	.B1(n36), 
	.B0(n942), 
	.A1(sboxw[18]), 
	.A0(n209));
   AOI222X1 U1273 (.Y(n1114), 
	.C1(n167), 
	.C0(n1553), 
	.B1(n37), 
	.B0(n359), 
	.A1(sboxw[2]), 
	.A0(n1557));
   OAI221XL U1274 (.Y(n1261), 
	.C0(n1268), 
	.B1(n318), 
	.B0(n1267), 
	.A1(n323), 
	.A0(sboxw[9]));
   AOI31X1 U1275 (.Y(n1268), 
	.B0(n1269), 
	.A2(n413), 
	.A1(n1511), 
	.A0(n50));
   NOR3BX1 U1276 (.Y(n1267), 
	.C(n571), 
	.B(n1270), 
	.AN(n316));
   OAI221XL U1277 (.Y(n1355), 
	.C0(n1368), 
	.B1(sboxw[13]), 
	.B0(n1367), 
	.A1(n318), 
	.A0(n1366));
   AOI222XL U1278 (.Y(n1366), 
	.C1(n1102), 
	.C0(n124), 
	.B1(n60), 
	.B0(n65), 
	.A1(n247), 
	.A0(n1507));
   AOI32XL U1279 (.Y(n1368), 
	.B1(sboxw[8]), 
	.B0(n286), 
	.A2(n291), 
	.A1(n24), 
	.A0(n290));
   AOI211XL U1280 (.Y(n1367), 
	.C0(n1370), 
	.B0(n1369), 
	.A1(n23), 
	.A0(n1503));
   OAI22X1 U1281 (.Y(n1460), 
	.B1(n1428), 
	.B0(sboxw[9]), 
	.A1(n156), 
	.A0(n1462));
   AOI211X1 U1282 (.Y(n1462), 
	.C0(n1301), 
	.B0(n1463), 
	.A1(n240), 
	.A0(n59));
   OAI21XL U1283 (.Y(n1463), 
	.B0(n1464), 
	.A1(n1311), 
	.A0(n55));
   AOI31XL U1284 (.Y(n1464), 
	.B0(n1341), 
	.A2(sboxw[12]), 
	.A1(n24), 
	.A0(n1278));
   AOI22X1 U1285 (.Y(n1017), 
	.B1(n33), 
	.B0(n211), 
	.A1(sboxw[18]), 
	.A0(n147));
   AOI22X1 U1286 (.Y(n434), 
	.B1(n34), 
	.B0(n1559), 
	.A1(sboxw[2]), 
	.A0(n166));
   OAI22X1 U1287 (.Y(new_sboxw[30]), 
	.B1(n1600), 
	.B0(n618), 
	.A1(n617), 
	.A0(sboxw[31]));
   AOI211X1 U1288 (.Y(n617), 
	.C0(n650), 
	.B0(n649), 
	.A1(n1598), 
	.A0(n648));
   AOI221X1 U1289 (.Y(n618), 
	.C0(n622), 
	.B1(n621), 
	.B0(n620), 
	.A1(n619), 
	.A0(sboxw[30]));
   OAI211X1 U1290 (.Y(n648), 
	.C0(n665), 
	.B0(n664), 
	.A1(n4), 
	.A0(n663));
   NOR2X1 U1291 (.Y(n988), 
	.B(sboxw[18]), 
	.A(n36));
   NOR2X1 U1292 (.Y(n405), 
	.B(sboxw[2]), 
	.A(n37));
   OAI221XL U1293 (.Y(n1306), 
	.C0(n1312), 
	.B1(n1308), 
	.B0(sboxw[9]), 
	.A1(n1311), 
	.A0(n55));
   AOI221XL U1294 (.Y(n1312), 
	.C0(n313), 
	.B1(n1517), 
	.B0(n1314), 
	.A1(n23), 
	.A0(n1313));
   AOI221X1 U1295 (.Y(n224), 
	.C0(n235), 
	.B1(n234), 
	.B0(n413), 
	.A1(n233), 
	.A0(n153));
   OAI221XL U1296 (.Y(n234), 
	.C0(n244), 
	.B1(n243), 
	.B0(n124), 
	.A1(n242), 
	.A0(sboxw[8]));
   OAI211XL U1297 (.Y(n233), 
	.C0(n249), 
	.B0(n248), 
	.A1(n247), 
	.A0(n246));
   AOI31X1 U1298 (.Y(n235), 
	.B0(n153), 
	.A2(n238), 
	.A1(n237), 
	.A0(n236));
   OAI211X1 U1299 (.Y(n879), 
	.C0(n888), 
	.B0(n887), 
	.A1(n881), 
	.A0(n138));
   AOI31X1 U1300 (.Y(n887), 
	.B0(n1567), 
	.A2(n577), 
	.A1(sboxw[28]), 
	.A0(n30));
   AOI222X1 U1301 (.Y(n888), 
	.C1(n136), 
	.C0(n1579), 
	.B1(n128), 
	.B0(n890), 
	.A1(n889), 
	.A0(n130));
   INVX1 U1302 (.Y(n1567), 
	.A(n655));
   OAI211X1 U1303 (.Y(n1228), 
	.C0(n1237), 
	.B0(n1236), 
	.A1(n1230), 
	.A0(n151));
   AOI31X1 U1304 (.Y(n1236), 
	.B0(n182), 
	.A2(n931), 
	.A1(sboxw[20]), 
	.A0(n29));
   AOI222X1 U1305 (.Y(n1237), 
	.C1(n146), 
	.C0(n179), 
	.B1(n142), 
	.B0(n1239), 
	.A1(n1238), 
	.A0(sboxw[21]));
   INVX1 U1306 (.Y(n182), 
	.A(n1009));
   OAI211X1 U1307 (.Y(n1472), 
	.C0(n1481), 
	.B0(n1480), 
	.A1(n1474), 
	.A0(n170));
   AOI31X1 U1308 (.Y(n1480), 
	.B0(n1529), 
	.A2(n348), 
	.A1(sboxw[4]), 
	.A0(n31));
   AOI222X1 U1309 (.Y(n1481), 
	.C1(n167), 
	.C0(n1526), 
	.B1(n160), 
	.B0(n1483), 
	.A1(n1482), 
	.A0(sboxw[5]));
   INVX1 U1310 (.Y(n1529), 
	.A(n426));
   OAI21XL U1311 (.Y(n995), 
	.B0(n151), 
	.A1(n203), 
	.A0(n187));
   OAI31X1 U1312 (.Y(n1440), 
	.B0(n1384), 
	.A2(n50), 
	.A1(sboxw[12]), 
	.A0(n1278));
   OAI22XL U1313 (.Y(n1302), 
	.B1(n125), 
	.B0(n254), 
	.A1(n12), 
	.A0(sboxw[9]));
   OAI221XL U1314 (.Y(n1456), 
	.C0(n1458), 
	.B1(sboxw[9]), 
	.B0(n17), 
	.A1(n124), 
	.A0(n1308));
   AOI211X1 U1315 (.Y(n1019), 
	.C0(n1022), 
	.B0(n1021), 
	.A1(n1020), 
	.A0(n931));
   OAI21XL U1316 (.Y(n1020), 
	.B0(sboxw[19]), 
	.A1(n36), 
	.A0(sboxw[20]));
   AOI21X1 U1317 (.Y(n1021), 
	.B0(n958), 
	.A1(n929), 
	.A0(n1023));
   NOR2X1 U1318 (.Y(n980), 
	.B(sboxw[20]), 
	.A(n1160));
   NOR2X1 U1319 (.Y(n397), 
	.B(sboxw[4]), 
	.A(n549));
   NAND2X1 U1320 (.Y(n314), 
	.B(n1515), 
	.A(sboxw[11]));
   OAI21XL U1321 (.Y(new_sboxw[28]), 
	.B0(n744), 
	.A1(n1600), 
	.A0(n743));
   AOI222X1 U1322 (.Y(n743), 
	.C1(n764), 
	.C0(n620), 
	.B1(n763), 
	.B0(n1595), 
	.A1(n762), 
	.A0(sboxw[30]));
   OAI2BB1X1 U1323 (.Y(n744), 
	.B0(n1600), 
	.A1N(n746), 
	.A0N(n745));
   OAI211X1 U1324 (.Y(n764), 
	.C0(n765), 
	.B0(n647), 
	.A1(n123), 
	.A0(n643));
   AOI31X1 U1325 (.Y(n785), 
	.B0(n557), 
	.A2(n788), 
	.A1(n787), 
	.A0(n786));
   NAND3X1 U1326 (.Y(n787), 
	.C(n1581), 
	.B(n730), 
	.A(sboxw[25]));
   AOI31X1 U1327 (.Y(n786), 
	.B0(n795), 
	.A2(n577), 
	.A1(sboxw[28]), 
	.A0(n137));
   AOI211X1 U1328 (.Y(n788), 
	.C0(n791), 
	.B0(n790), 
	.A1(n26), 
	.A0(n789));
   AOI31X1 U1329 (.Y(n1134), 
	.B0(n911), 
	.A2(n1137), 
	.A1(n1136), 
	.A0(n1135));
   NAND3X1 U1330 (.Y(n1136), 
	.C(n181), 
	.B(n1051), 
	.A(sboxw[17]));
   AOI31X1 U1331 (.Y(n1135), 
	.B0(n1144), 
	.A2(n931), 
	.A1(sboxw[20]), 
	.A0(n150));
   AOI211X1 U1332 (.Y(n1137), 
	.C0(n1140), 
	.B0(n1139), 
	.A1(n27), 
	.A0(n1138));
   AOI31X1 U1333 (.Y(n523), 
	.B0(n328), 
	.A2(n526), 
	.A1(n525), 
	.A0(n524));
   NAND3X1 U1334 (.Y(n525), 
	.C(n1528), 
	.B(n468), 
	.A(sboxw[1]));
   AOI31X1 U1335 (.Y(n524), 
	.B0(n533), 
	.A2(n348), 
	.A1(sboxw[4]), 
	.A0(n168));
   AOI211X1 U1336 (.Y(n526), 
	.C0(n529), 
	.B0(n528), 
	.A1(n28), 
	.A0(n527));
   NAND2X1 U1337 (.Y(n1394), 
	.B(n1511), 
	.A(sboxw[10]));
   AOI32XL U1338 (.Y(n225), 
	.B1(n228), 
	.B0(n219), 
	.A2(n227), 
	.A1(n24), 
	.A0(sboxw[14]));
   OAI221XL U1339 (.Y(n228), 
	.C0(n231), 
	.B1(n24), 
	.B0(n230), 
	.A1(n12), 
	.A0(n65));
   AOI211X1 U1340 (.Y(n231), 
	.C0(n925), 
	.B0(n232), 
	.A1(n59), 
	.A0(n127));
   OAI211XL U1341 (.Y(n1465), 
	.C0(n1458), 
	.B0(n1334), 
	.A1(n12), 
	.A0(sboxw[9]));
   NAND2X1 U1342 (.Y(n1334), 
	.B(sboxw[8]), 
	.A(n1506));
   NOR2X1 U1343 (.Y(n1314), 
	.B(sboxw[12]), 
	.A(n1510));
   NAND2X1 U1344 (.Y(n1289), 
	.B(sboxw[9]), 
	.A(n59));
   AOI31X1 U1345 (.Y(n1431), 
	.B0(n1435), 
	.A2(n1434), 
	.A1(n1433), 
	.A0(n1432));
   AOI22X1 U1346 (.Y(n1432), 
	.B1(n1503), 
	.B0(n127), 
	.A1(sboxw[8]), 
	.A0(n739));
   AOI222X1 U1347 (.Y(n1434), 
	.C1(n50), 
	.C0(n1506), 
	.B1(n1517), 
	.B0(n59), 
	.A1(n60), 
	.A0(n1336));
   AOI21X1 U1348 (.Y(n1433), 
	.B0(n1060), 
	.A1(n635), 
	.A0(n65));
   AOI31X1 U1349 (.Y(n1273), 
	.B0(n223), 
	.A2(n1276), 
	.A1(n1275), 
	.A0(n1274));
   AOI31XL U1350 (.Y(n1274), 
	.B0(n263), 
	.A2(n65), 
	.A1(n242), 
	.A0(sboxw[10]));
   AOI22X1 U1351 (.Y(n1276), 
	.B1(n55), 
	.B0(n739), 
	.A1(n1277), 
	.A0(sboxw[8]));
   NAND3X1 U1352 (.Y(n1275), 
	.C(sboxw[12]), 
	.B(n125), 
	.A(n1278));
   AOI22XL U1353 (.Y(n1458), 
	.B1(n59), 
	.B0(n23), 
	.A1(sboxw[9]), 
	.A0(n1061));
   AOI31X1 U1354 (.Y(n1272), 
	.B0(sboxw[14]), 
	.A2(n1281), 
	.A1(n1280), 
	.A0(n1279));
   AOI31X1 U1355 (.Y(n1280), 
	.B0(n1286), 
	.A2(n291), 
	.A1(n1511), 
	.A0(n126));
   AOI2BB2X1 U1356 (.Y(n1279), 
	.B1(n1507), 
	.B0(n1287), 
	.A1N(n65), 
	.A0N(n1288));
   AOI221X1 U1357 (.Y(n1281), 
	.C0(n1282), 
	.B1(n25), 
	.B0(n227), 
	.A1(sboxw[9]), 
	.A0(n1503));
   AOI31X1 U1358 (.Y(n560), 
	.B0(sboxw[30]), 
	.A2(n570), 
	.A1(n569), 
	.A0(n568));
   AOI2BB2X1 U1359 (.Y(n568), 
	.B1(n1593), 
	.B0(n579), 
	.A1N(n30), 
	.A0N(n580));
   AOI31X1 U1360 (.Y(n569), 
	.B0(n578), 
	.A2(n577), 
	.A1(n1592), 
	.A0(n576));
   AOI221X1 U1361 (.Y(n570), 
	.C0(n572), 
	.B1(n10), 
	.B0(n1577), 
	.A1(n135), 
	.A0(n1574));
   AOI31X1 U1362 (.Y(n1282), 
	.B0(sboxw[13]), 
	.A2(n1285), 
	.A1(n1284), 
	.A0(n1283));
   AOI21X1 U1363 (.Y(n1285), 
	.B0(n1270), 
	.A1(n1061), 
	.A0(sboxw[9]));
   AOI21X1 U1364 (.Y(n742), 
	.B0(n599), 
	.A1(n734), 
	.A0(n598));
   AOI31X1 U1365 (.Y(n1056), 
	.B0(n1063), 
	.A2(n185), 
	.A1(n970), 
	.A0(sboxw[20]));
   AOI21X1 U1366 (.Y(n1063), 
	.B0(n953), 
	.A1(n1055), 
	.A0(n952));
   AOI31X1 U1367 (.Y(n473), 
	.B0(n480), 
	.A2(n1532), 
	.A1(n387), 
	.A0(sboxw[4]));
   AOI21X1 U1368 (.Y(n480), 
	.B0(n370), 
	.A1(n472), 
	.A0(n369));
   AOI31XL U1369 (.Y(n1372), 
	.B0(n1378), 
	.A2(n413), 
	.A1(n247), 
	.A0(sboxw[12]));
   AOI21X1 U1370 (.Y(n1378), 
	.B0(n318), 
	.A1(n324), 
	.A0(n316));
   OAI22X1 U1371 (.Y(n649), 
	.B1(n657), 
	.B0(n656), 
	.A1(n655), 
	.A0(n1598));
   AOI211X1 U1372 (.Y(n656), 
	.C0(n659), 
	.B0(n658), 
	.A1(n138), 
	.A0(n1576));
   OAI21XL U1373 (.Y(n659), 
	.B0(n661), 
	.A1(n660), 
	.A0(n123));
   OAI222XL U1374 (.Y(n658), 
	.C1(n662), 
	.C0(sboxw[28]), 
	.B1(n643), 
	.B0(n135), 
	.A1(n11), 
	.A0(n22));
   OAI22X1 U1375 (.Y(n1003), 
	.B1(n1011), 
	.B0(n1010), 
	.A1(n1009), 
	.A0(n174));
   AOI211X1 U1376 (.Y(n1010), 
	.C0(n1013), 
	.B0(n1012), 
	.A1(n151), 
	.A0(n202));
   OAI21XL U1377 (.Y(n1013), 
	.B0(n1015), 
	.A1(n1014), 
	.A0(n120));
   OAI222XL U1378 (.Y(n1012), 
	.C1(n1016), 
	.C0(sboxw[20]), 
	.B1(n997), 
	.B0(n147), 
	.A1(n8), 
	.A0(n999));
   OAI22X1 U1379 (.Y(n420), 
	.B1(n428), 
	.B0(n427), 
	.A1(n426), 
	.A0(n1521));
   AOI211X1 U1380 (.Y(n427), 
	.C0(n430), 
	.B0(n429), 
	.A1(n170), 
	.A0(n1550));
   OAI21XL U1381 (.Y(n430), 
	.B0(n432), 
	.A1(n431), 
	.A0(n117));
   OAI222XL U1382 (.Y(n429), 
	.C1(n433), 
	.C0(sboxw[4]), 
	.B1(n414), 
	.B0(sboxw[1]), 
	.A1(n7), 
	.A0(n416));
   NAND2X1 U1383 (.Y(n298), 
	.B(sboxw[9]), 
	.A(n1502));
   NAND2X1 U1384 (.Y(n669), 
	.B(sboxw[27]), 
	.A(n30));
   NAND2X1 U1385 (.Y(n1023), 
	.B(sboxw[19]), 
	.A(n29));
   NAND2X1 U1386 (.Y(n440), 
	.B(sboxw[3]), 
	.A(n31));
   NAND2X1 U1387 (.Y(n1428), 
	.B(sboxw[11]), 
	.A(n291));
   OAI22X1 U1388 (.Y(n1324), 
	.B1(n1330), 
	.B0(n1329), 
	.A1(n304), 
	.A0(n217));
   AOI211X1 U1389 (.Y(n1329), 
	.C0(n902), 
	.B0(n1332), 
	.A1(n1251), 
	.A0(n1331));
   OAI221XL U1390 (.Y(n1332), 
	.C0(n1334), 
	.B1(n1311), 
	.B0(sboxw[8]), 
	.A1(n1333), 
	.A0(n24));
   INVX1 U1391 (.Y(n902), 
	.A(n315));
   AOI31X1 U1392 (.Y(n561), 
	.B0(n565), 
	.A2(n564), 
	.A1(n563), 
	.A0(n562));
   NAND3X1 U1393 (.Y(n563), 
	.C(n51), 
	.B(sboxw[26]), 
	.A(n30));
   AOI31X1 U1394 (.Y(n562), 
	.B0(n567), 
	.A2(n26), 
	.A1(n1572), 
	.A0(sboxw[28]));
   AOI22X1 U1395 (.Y(n564), 
	.B1(n32), 
	.B0(n1575), 
	.A1(n566), 
	.A0(n137));
   AOI31X1 U1396 (.Y(n915), 
	.B0(n919), 
	.A2(n918), 
	.A1(n917), 
	.A0(n916));
   NAND3X1 U1397 (.Y(n917), 
	.C(n52), 
	.B(sboxw[18]), 
	.A(n29));
   AOI31X1 U1398 (.Y(n916), 
	.B0(n921), 
	.A2(n27), 
	.A1(n206), 
	.A0(sboxw[20]));
   AOI22X1 U1399 (.Y(n918), 
	.B1(n33), 
	.B0(n190), 
	.A1(n920), 
	.A0(n150));
   AOI31X1 U1400 (.Y(n332), 
	.B0(n336), 
	.A2(n335), 
	.A1(n334), 
	.A0(n333));
   NAND3X1 U1401 (.Y(n334), 
	.C(n53), 
	.B(sboxw[2]), 
	.A(n31));
   AOI31X1 U1402 (.Y(n333), 
	.B0(n338), 
	.A2(n28), 
	.A1(n1554), 
	.A0(sboxw[4]));
   AOI22X1 U1403 (.Y(n335), 
	.B1(n34), 
	.B0(n1538), 
	.A1(n337), 
	.A0(n168));
   AOI22X1 U1404 (.Y(n745), 
	.B1(n752), 
	.B0(sboxw[30]), 
	.A1(n751), 
	.A0(n620));
   OAI221XL U1405 (.Y(n751), 
	.C0(n761), 
	.B1(n4), 
	.B0(n30), 
	.A1(n642), 
	.A0(n26));
   OAI222XL U1406 (.Y(n752), 
	.C1(n129), 
	.C0(n755), 
	.B1(n599), 
	.B0(n754), 
	.A1(n753), 
	.A0(n130));
   AOI211X1 U1407 (.Y(n761), 
	.C0(n589), 
	.B0(n1586), 
	.A1(n135), 
	.A0(n629));
   AOI22X1 U1408 (.Y(n483), 
	.B1(n490), 
	.B0(sboxw[6]), 
	.A1(n489), 
	.A0(n391));
   OAI221XL U1409 (.Y(n489), 
	.C0(n499), 
	.B1(n16), 
	.B0(n31), 
	.A1(n9), 
	.A0(n28));
   OAI222XL U1410 (.Y(n490), 
	.C1(n161), 
	.C0(n493), 
	.B1(n370), 
	.B0(n492), 
	.A1(n491), 
	.A0(n159));
   AOI211X1 U1411 (.Y(n499), 
	.C0(n360), 
	.B0(n62), 
	.A1(sboxw[1]), 
	.A0(n400));
   AOI22X1 U1412 (.Y(n1381), 
	.B1(n1388), 
	.B0(sboxw[14]), 
	.A1(n1387), 
	.A0(n215));
   OAI221XL U1413 (.Y(n1387), 
	.C0(n1395), 
	.B1(n13), 
	.B0(n65), 
	.A1(n240), 
	.A0(n243));
   OAI222XL U1414 (.Y(n1388), 
	.C1(n156), 
	.C0(n1391), 
	.B1(n318), 
	.B0(n1390), 
	.A1(n1389), 
	.A0(n153));
   AOI211X1 U1415 (.Y(n1395), 
	.C0(n1266), 
	.B0(n59), 
	.A1(sboxw[9]), 
	.A0(n1313));
   AOI22X1 U1416 (.Y(n1018), 
	.B1(n142), 
	.B0(n1025), 
	.A1(n1024), 
	.A0(sboxw[21]));
   OAI21XL U1417 (.Y(n1024), 
	.B0(n948), 
	.A1(n1026), 
	.A0(n147));
   OAI22X1 U1418 (.Y(n1025), 
	.B1(n999), 
	.B0(n1017), 
	.A1(n33), 
	.A0(sboxw[19]));
   AOI22X1 U1419 (.Y(n435), 
	.B1(n161), 
	.B0(n442), 
	.A1(n441), 
	.A0(n159));
   OAI21XL U1420 (.Y(n441), 
	.B0(n365), 
	.A1(n443), 
	.A0(n166));
   OAI22X1 U1421 (.Y(n442), 
	.B1(n416), 
	.B0(n434), 
	.A1(n34), 
	.A0(sboxw[3]));
   AND2X2 U1422 (.Y(n54), 
	.B(n1517), 
	.A(sboxw[9]));
   NAND4X1 U1424 (.Y(n1383), 
	.D(n1386), 
	.C(n1385), 
	.B(n1284), 
	.A(n1384));
   NAND3X1 U1425 (.Y(n1385), 
	.C(sboxw[10]), 
	.B(n23), 
	.A(n290));
   AOI222X1 U1426 (.Y(n1386), 
	.C1(n25), 
	.C0(n739), 
	.B1(n50), 
	.B0(n1314), 
	.A1(n1503), 
	.A0(n55));
   INVX1 U1428 (.Y(n1516), 
	.A(sboxw[9]));
   NAND4X1 U1429 (.Y(n1412), 
	.D(n1423), 
	.C(n1422), 
	.B(n1421), 
	.A(n1420));
   NAND3X1 U1430 (.Y(n1423), 
	.C(n49), 
	.B(n290), 
	.A(sboxw[9]));
   AOI22X1 U1431 (.Y(n1420), 
	.B1(n125), 
	.B0(n477), 
	.A1(n156), 
	.A0(n1427));
   AOI31X1 U1432 (.Y(n1422), 
	.B0(n229), 
	.A2(n291), 
	.A1(sboxw[12]), 
	.A0(sboxw[8]));
   NAND4X1 U1433 (.Y(n1271), 
	.D(n1292), 
	.C(n1291), 
	.B(n1290), 
	.A(n1289));
   AOI221XL U1434 (.Y(n1292), 
	.C0(n277), 
	.B1(n25), 
	.B0(n1506), 
	.A1(n24), 
	.A0(n1503));
   AOI21X1 U1435 (.Y(n1291), 
	.B0(n1266), 
	.A1(sboxw[8]), 
	.A0(n239));
   OAI2BB2X1 U1436 (.Y(n1430), 
	.B1(n1330), 
	.B0(n1436), 
	.A1N(n1437), 
	.A0N(n218));
   NAND4X1 U1437 (.Y(n1437), 
	.D(n1438), 
	.C(n1326), 
	.B(n230), 
	.A(n1401));
   AOI211X1 U1438 (.Y(n1436), 
	.C0(n1440), 
	.B0(n1439), 
	.A1(sboxw[10]), 
	.A0(n55));
   AOI222X1 U1439 (.Y(n1438), 
	.C1(n1512), 
	.C0(n55), 
	.B1(n1517), 
	.B0(n301), 
	.A1(n1102), 
	.A0(n1336));
   NAND4BXL U1440 (.Y(n819), 
	.D(n833), 
	.C(n832), 
	.B(n661), 
	.AN(n628));
   AOI22X1 U1441 (.Y(n832), 
	.B1(sboxw[26]), 
	.B0(n1568), 
	.A1(n26), 
	.A0(n758));
   AOI222X1 U1442 (.Y(n833), 
	.C1(n123), 
	.C0(n1582), 
	.B1(n136), 
	.B0(n1576), 
	.A1(n11), 
	.A0(n1591));
   NAND4BXL U1443 (.Y(n1168), 
	.D(n1182), 
	.C(n1181), 
	.B(n1015), 
	.AN(n982));
   AOI22X1 U1444 (.Y(n1181), 
	.B1(sboxw[18]), 
	.B0(n209), 
	.A1(n27), 
	.A0(n1079));
   AOI222X1 U1445 (.Y(n1182), 
	.C1(n120), 
	.C0(n187), 
	.B1(n146), 
	.B0(n202), 
	.A1(n8), 
	.A0(n196));
   NAND4BXL U1446 (.Y(n676), 
	.D(n690), 
	.C(n689), 
	.B(n432), 
	.AN(n399));
   AOI22X1 U1447 (.Y(n689), 
	.B1(sboxw[2]), 
	.B0(n1557), 
	.A1(n28), 
	.A0(n496));
   AOI222X1 U1448 (.Y(n690), 
	.C1(n117), 
	.C0(n1534), 
	.B1(n167), 
	.B0(n1550), 
	.A1(n7), 
	.A0(n1544));
   NAND4BXL U1449 (.Y(n256), 
	.D(n266), 
	.C(n265), 
	.B(n264), 
	.AN(n263));
   AOI22X1 U1450 (.Y(n265), 
	.B1(n1495), 
	.B0(sboxw[8]), 
	.A1(n25), 
	.A0(n252));
   AOI222X1 U1451 (.Y(n266), 
	.C1(n59), 
	.C0(n124), 
	.B1(n240), 
	.B0(n1503), 
	.A1(n50), 
	.A0(n1502));
   OAI21XL U1452 (.Y(n962), 
	.B0(n964), 
	.A1(n963), 
	.A0(sboxw[20]));
   AOI22X1 U1453 (.Y(n963), 
	.B1(n181), 
	.B0(n38), 
	.A1(n119), 
	.A0(n931));
   OAI21XL U1454 (.Y(n379), 
	.B0(n381), 
	.A1(n380), 
	.A0(sboxw[4]));
   AOI22X1 U1455 (.Y(n380), 
	.B1(n1528), 
	.B0(n39), 
	.A1(n116), 
	.A0(n348));
   NAND4X1 U1456 (.Y(n763), 
	.D(n771), 
	.C(n770), 
	.B(n769), 
	.A(n768));
   NAND3X1 U1457 (.Y(n770), 
	.C(n51), 
	.B(n11), 
	.A(sboxw[26]));
   AOI222X1 U1458 (.Y(n771), 
	.C1(n35), 
	.C0(n1575), 
	.B1(n135), 
	.B0(n772), 
	.A1(n10), 
	.A0(n1586));
   NAND4X1 U1459 (.Y(n501), 
	.D(n509), 
	.C(n508), 
	.B(n507), 
	.A(n506));
   NAND3X1 U1460 (.Y(n508), 
	.C(n53), 
	.B(n115), 
	.A(sboxw[2]));
   AOI222X1 U1461 (.Y(n509), 
	.C1(n37), 
	.C0(n1538), 
	.B1(n166), 
	.B0(n510), 
	.A1(n116), 
	.A0(n62));
   NAND4X1 U1462 (.Y(n1397), 
	.D(n1403), 
	.C(n1402), 
	.B(n249), 
	.A(n1401));
   NAND3X1 U1463 (.Y(n1402), 
	.C(n645), 
	.B(n23), 
	.A(sboxw[10]));
   AOI222X1 U1464 (.Y(n1403), 
	.C1(n124), 
	.C0(n739), 
	.B1(sboxw[9]), 
	.B0(n1512), 
	.A1(n25), 
	.A0(n59));
   NAND4X1 U1465 (.Y(n1413), 
	.D(n1416), 
	.C(n1415), 
	.B(n1414), 
	.A(n1296));
   AOI22X1 U1466 (.Y(n1415), 
	.B1(n58), 
	.B0(n1287), 
	.A1(n55), 
	.A0(n1335));
   AOI211X1 U1467 (.Y(n1416), 
	.C0(n1364), 
	.B0(n1417), 
	.A1(sboxw[9]), 
	.A0(n477));
   AOI21X1 U1468 (.Y(n1417), 
	.B0(sboxw[13]), 
	.A1(n1419), 
	.A0(n1418));
   OAI21XL U1469 (.Y(n641), 
	.B0(n139), 
	.A1(n66), 
	.A0(n1582));
   OAI21XL U1470 (.Y(n412), 
	.B0(n169), 
	.A1(n1551), 
	.A0(n1534));
   AND2X2 U1471 (.Y(n55), 
	.B(n1516), 
	.A(sboxw[8]));
   AOI21X1 U1472 (.Y(n934), 
	.B0(n935), 
	.A1(n181), 
	.A0(sboxw[20]));
   AOI21X1 U1473 (.Y(n351), 
	.B0(n352), 
	.A1(n1528), 
	.A0(sboxw[4]));
   AOI21X1 U1474 (.Y(n1288), 
	.B0(n271), 
	.A1(n49), 
	.A0(sboxw[12]));
   AND2X2 U1475 (.Y(n56), 
	.B(sboxw[19]), 
	.A(sboxw[20]));
   INVX1 U1476 (.Y(n999), 
	.A(n56));
   AND2X2 U1477 (.Y(n57), 
	.B(sboxw[3]), 
	.A(sboxw[4]));
   INVX1 U1478 (.Y(n416), 
	.A(n57));
   AND2X2 U1479 (.Y(n1269), 
	.B(sboxw[9]), 
	.A(n274));
   INVX1 U1480 (.Y(n1517), 
	.A(sboxw[8]));
   INVX1 U1481 (.Y(n1515), 
	.A(sboxw[10]));
   INVX1 U1482 (.Y(n211), 
	.A(sboxw[18]));
   INVX1 U1483 (.Y(n1559), 
	.A(sboxw[2]));
   AND2X2 U1484 (.Y(n58), 
	.B(n1251), 
	.A(sboxw[11]));
   INVX1 U1485 (.Y(n243), 
	.A(n58));
   AND2X2 U1486 (.Y(n59), 
	.B(sboxw[10]), 
	.A(n58));
   INVX1 U1487 (.Y(n254), 
	.A(n59));
   AND2X2 U1488 (.Y(n60), 
	.B(n1511), 
	.A(sboxw[12]));
   INVX1 U1489 (.Y(n242), 
	.A(n60));
   INVX1 U1490 (.Y(n1592), 
	.A(sboxw[27]));
   INVX1 U1491 (.Y(n207), 
	.A(sboxw[19]));
   INVX1 U1492 (.Y(n1555), 
	.A(sboxw[3]));
   AND2X2 U1493 (.Y(n61), 
	.B(n64), 
	.A(sboxw[18]));
   INVX1 U1494 (.Y(n1026), 
	.A(n61));
   AND2X2 U1495 (.Y(n62), 
	.B(n1536), 
	.A(sboxw[2]));
   INVX1 U1496 (.Y(n443), 
	.A(n62));
   INVX1 U1497 (.Y(n1511), 
	.A(sboxw[11]));
   AND2X2 U1498 (.Y(n63), 
	.B(n1594), 
	.A(sboxw[27]));
   INVX1 U1499 (.Y(n642), 
	.A(n63));
   AND2X2 U1500 (.Y(n64), 
	.B(n197), 
	.A(sboxw[19]));
   INVX1 U1501 (.Y(n996), 
	.A(n64));
   INVX1 U1502 (.Y(n138), 
	.A(sboxw[24]));
   INVX1 U1505 (.Y(n169), 
	.A(sboxw[0]));
   INVX1 U1506 (.Y(n146), 
	.A(sboxw[17]));
   INVX1 U1509 (.Y(n159), 
	.A(n160));
   INVX1 U1510 (.Y(n174), 
	.A(sboxw[22]));
   INVX1 U1511 (.Y(n1521), 
	.A(sboxw[6]));
   NOR2X1 U1512 (.Y(n758), 
	.B(sboxw[27]), 
	.A(n1583));
   NOR2X1 U1513 (.Y(n974), 
	.B(sboxw[22]), 
	.A(n142));
   NOR2X1 U1514 (.Y(n391), 
	.B(sboxw[6]), 
	.A(n161));
   AOI22X1 U1515 (.Y(n1336), 
	.B1(n55), 
	.B0(n1515), 
	.A1(sboxw[9]), 
	.A0(sboxw[10]));
   NOR2X1 U1516 (.Y(n239), 
	.B(sboxw[11]), 
	.A(sboxw[10]));
   NOR2X1 U1517 (.Y(n942), 
	.B(sboxw[19]), 
	.A(sboxw[18]));
   NOR2X1 U1518 (.Y(n359), 
	.B(sboxw[3]), 
	.A(sboxw[2]));
   OAI222XL U1519 (.Y(n1439), 
	.C1(n12), 
	.C0(n127), 
	.B1(n1517), 
	.B0(n1374), 
	.A1(n1308), 
	.A0(sboxw[8]));
   AOI222X1 U1520 (.Y(n238), 
	.C1(n1516), 
	.C0(n1508), 
	.B1(n124), 
	.B0(n239), 
	.A1(sboxw[10]), 
	.A0(n1513));
   NOR2X1 U1521 (.Y(n772), 
	.B(sboxw[26]), 
	.A(n1592));
   NOR2X1 U1522 (.Y(n1093), 
	.B(sboxw[18]), 
	.A(n207));
   NOR2X1 U1523 (.Y(n510), 
	.B(sboxw[2]), 
	.A(n1555));
   NOR2X1 U1524 (.Y(n312), 
	.B(sboxw[10]), 
	.A(n1251));
   AOI22X1 U1525 (.Y(n663), 
	.B1(n32), 
	.B0(n1583), 
	.A1(sboxw[26]), 
	.A0(n135));
   NAND2X1 U1526 (.Y(n1333), 
	.B(sboxw[10]), 
	.A(sboxw[12]));
   NOR2X1 U1527 (.Y(n301), 
	.B(sboxw[12]), 
	.A(n1515));
   AOI22X1 U1528 (.Y(n1321), 
	.B1(n55), 
	.B0(sboxw[10]), 
	.A1(n1515), 
	.A0(n1517));
   NOR2X1 U1529 (.Y(n780), 
	.B(sboxw[28]), 
	.A(n1583));
   NOR2X1 U1530 (.Y(n1101), 
	.B(sboxw[20]), 
	.A(n211));
   NOR2X1 U1531 (.Y(n518), 
	.B(sboxw[4]), 
	.A(n1559));
   NOR2X1 U1532 (.Y(n634), 
	.B(sboxw[26]), 
	.A(n35));
   OAI221XL U1533 (.Y(n1351), 
	.C0(sboxw[11]), 
	.B1(sboxw[12]), 
	.B0(sboxw[8]), 
	.A1(n1251), 
	.A0(n124));
   OAI221XL U1534 (.Y(n711), 
	.C0(sboxw[27]), 
	.B1(sboxw[24]), 
	.B0(sboxw[28]), 
	.A1(n1594), 
	.A0(n35));
   OAI221XL U1535 (.Y(n1032), 
	.C0(sboxw[19]), 
	.B1(sboxw[16]), 
	.B0(sboxw[20]), 
	.A1(n197), 
	.A0(n36));
   OAI221XL U1536 (.Y(n449), 
	.C0(sboxw[3]), 
	.B1(sboxw[0]), 
	.B0(sboxw[4]), 
	.A1(n1545), 
	.A0(n37));
   NOR2X1 U1537 (.Y(n302), 
	.B(sboxw[10]), 
	.A(n124));
   AOI211X1 U1538 (.Y(n665), 
	.C0(n668), 
	.B0(n667), 
	.A1(n666), 
	.A0(n577));
   OAI21XL U1539 (.Y(n666), 
	.B0(sboxw[27]), 
	.A1(n35), 
	.A0(sboxw[28]));
   AOI21X1 U1540 (.Y(n667), 
	.B0(n604), 
	.A1(n575), 
	.A0(n669));
   AOI211X1 U1541 (.Y(n436), 
	.C0(n439), 
	.B0(n438), 
	.A1(n437), 
	.A0(n348));
   OAI21XL U1542 (.Y(n437), 
	.B0(sboxw[3]), 
	.A1(n37), 
	.A0(sboxw[4]));
   AOI21X1 U1543 (.Y(n438), 
	.B0(n375), 
	.A1(n346), 
	.A0(n440));
   NOR2X1 U1544 (.Y(n626), 
	.B(sboxw[28]), 
	.A(n811));
   OAI211X1 U1545 (.Y(n1085), 
	.C0(n1086), 
	.B0(n1001), 
	.A1(n120), 
	.A0(n997));
   AOI21X1 U1546 (.Y(n1086), 
	.B0(n1087), 
	.A1(n33), 
	.A0(n187));
   OAI211X1 U1547 (.Y(n502), 
	.C0(n503), 
	.B0(n418), 
	.A1(n117), 
	.A0(n414));
   AOI21X1 U1548 (.Y(n503), 
	.B0(n504), 
	.A1(n34), 
	.A0(n1534));
   NAND2X1 U1549 (.Y(n565), 
	.B(n129), 
	.A(sboxw[30]));
   NAND2X1 U1550 (.Y(n919), 
	.B(n142), 
	.A(sboxw[22]));
   NAND2X1 U1551 (.Y(n336), 
	.B(n161), 
	.A(sboxw[6]));
   NAND2X1 U1552 (.Y(n223), 
	.B(sboxw[13]), 
	.A(sboxw[14]));
   OAI22X1 U1553 (.Y(n1344), 
	.B1(n230), 
	.B0(n1336), 
	.A1(n55), 
	.A0(sboxw[11]));
   AOI31X1 U1554 (.Y(n293), 
	.B0(n342), 
	.A2(n291), 
	.A1(sboxw[12]), 
	.A0(n65));
   INVX1 U1555 (.Y(n342), 
	.A(n304));
   AOI22XL U1556 (.Y(n277), 
	.B1(sboxw[10]), 
	.B0(n24), 
	.A1(n247), 
	.A0(n1515));
   NAND3X1 U1557 (.Y(n768), 
	.C(n30), 
	.B(n1583), 
	.A(sboxw[28]));
   NAND3X1 U1558 (.Y(n1089), 
	.C(n29), 
	.B(n211), 
	.A(sboxw[20]));
   NAND3X1 U1559 (.Y(n506), 
	.C(n31), 
	.B(n1559), 
	.A(sboxw[4]));
   NAND2X1 U1560 (.Y(n324), 
	.B(n58), 
	.A(sboxw[8]));
   NAND2X1 U1561 (.Y(n1330), 
	.B(n153), 
	.A(sboxw[14]));
   NAND2X1 U1562 (.Y(n1014), 
	.B(sboxw[20]), 
	.A(sboxw[18]));
   NAND2X1 U1563 (.Y(n431), 
	.B(sboxw[4]), 
	.A(sboxw[2]));
   NOR2X1 U1564 (.Y(n982), 
	.B(sboxw[18]), 
	.A(n6));
   NOR2X1 U1565 (.Y(n399), 
	.B(sboxw[2]), 
	.A(n5));
   OAI21XL U1566 (.Y(n1343), 
	.B0(n258), 
	.A1(n254), 
	.A0(sboxw[9]));
   AOI22X1 U1567 (.Y(n244), 
	.B1(n1507), 
	.B0(sboxw[8]), 
	.A1(n25), 
	.A0(n1102));
   AND2X2 U1568 (.Y(n65), 
	.B(sboxw[9]), 
	.A(sboxw[8]));
   AOI22X1 U1570 (.Y(n664), 
	.B1(n129), 
	.B0(n671), 
	.A1(n670), 
	.A0(n130));
   OAI21XL U1571 (.Y(n670), 
	.B0(n594), 
	.A1(n14), 
	.A0(n135));
   OAI22X1 U1572 (.Y(n671), 
	.B1(n22), 
	.B0(n663), 
	.A1(n32), 
	.A0(sboxw[27]));
   OAI21XL U1573 (.Y(n1294), 
	.B0(n1296), 
	.A1(n1295), 
	.A0(sboxw[12]));
   AOI22X1 U1574 (.Y(n1295), 
	.B1(n50), 
	.B0(n49), 
	.A1(n25), 
	.A0(n291));
   OAI21XL U1575 (.Y(n608), 
	.B0(n610), 
	.A1(n609), 
	.A0(sboxw[28]));
   AOI22X1 U1576 (.Y(n609), 
	.B1(n1581), 
	.B0(n40), 
	.A1(n122), 
	.A0(n577));
   NAND2X1 U1577 (.Y(n1361), 
	.B(sboxw[11]), 
	.A(n65));
   OAI21XL U1578 (.Y(n1339), 
	.B0(sboxw[11]), 
	.A1(n54), 
	.A0(sboxw[12]));
   AOI21X1 U1579 (.Y(n765), 
	.B0(n766), 
	.A1(n32), 
	.A0(n1582));
   AOI21X1 U1580 (.Y(n580), 
	.B0(n581), 
	.A1(n1581), 
	.A0(sboxw[28]));
   AND2X2 U1581 (.Y(n66), 
	.B(n1590), 
	.A(sboxw[26]));
   INVX1 U1582 (.Y(n740), 
	.A(n66));
   INVX1 U1583 (.Y(n1583), 
	.A(sboxw[26]));
   AOI211X1 U1584 (.Y(n222), 
	.C0(n251), 
	.B0(n250), 
	.A1(n1503), 
	.A0(n124));
   OAI222XL U1585 (.Y(n250), 
	.C1(n24), 
	.C0(n243), 
	.B1(n254), 
	.B0(sboxw[8]), 
	.A1(n12), 
	.A0(n50));
   OAI2BB1X1 U1586 (.Y(n251), 
	.B0(n253), 
	.A1N(n127), 
	.A0N(n252));
   OAI21XL U1587 (.Y(n253), 
	.B0(sboxw[8]), 
	.A1(n1061), 
	.A0(n1495));
   AND2X2 U1588 (.Y(n67), 
	.B(n1593), 
	.A(sboxw[26]));
   INVX1 U1589 (.Y(n781), 
	.A(n67));
   INVX1 U1591 (.Y(n1598), 
	.A(sboxw[30]));
   NOR2X1 U1592 (.Y(n620), 
	.B(sboxw[30]), 
	.A(n129));
   NOR2X1 U1593 (.Y(n588), 
	.B(sboxw[27]), 
	.A(sboxw[26]));
   OAI22X1 U1594 (.Y(n275), 
	.B1(n242), 
	.B0(sboxw[9]), 
	.A1(n1516), 
	.A0(n1511));
   NAND2X1 U1595 (.Y(n557), 
	.B(n1598), 
	.A(sboxw[31]));
   NAND2X1 U1596 (.Y(n911), 
	.B(n174), 
	.A(sboxw[23]));
   NAND2X1 U1597 (.Y(n328), 
	.B(n1521), 
	.A(sboxw[7]));
   AOI22X1 U1598 (.Y(n297), 
	.B1(sboxw[10]), 
	.B0(n24), 
	.A1(sboxw[8]), 
	.A0(n1515));
   NAND2X1 U1599 (.Y(n660), 
	.B(sboxw[28]), 
	.A(sboxw[26]));
   NAND2X1 U1600 (.Y(n657), 
	.B(n130), 
	.A(sboxw[30]));
   NAND2X1 U1601 (.Y(n1011), 
	.B(n143), 
	.A(sboxw[22]));
   NAND2X1 U1602 (.Y(n428), 
	.B(n159), 
	.A(sboxw[6]));
   NAND2X1 U1603 (.Y(n1346), 
	.B(n217), 
	.A(sboxw[15]));
   NOR2X1 U1604 (.Y(n628), 
	.B(sboxw[26]), 
	.A(n10));
   NAND2X1 U1605 (.Y(n1326), 
	.B(sboxw[8]), 
	.A(n1508));
   INVX1 U1606 (.Y(n217), 
	.A(sboxw[14]));
   INVX1 U1607 (.Y(n1600), 
	.A(sboxw[31]));
   INVX1 U1608 (.Y(n212), 
	.A(sboxw[15]));
   INVX1 U1609 (.Y(n171), 
	.A(sboxw[23]));
   INVX1 U1610 (.Y(n1518), 
	.A(sboxw[7]));
   NAND2X1 U1611 (.Y(n1258), 
	.B(sboxw[14]), 
	.A(sboxw[15]));
   NAND2X1 U1612 (.Y(n555), 
	.B(sboxw[31]), 
	.A(sboxw[30]));
   NAND2X1 U1613 (.Y(n909), 
	.B(sboxw[23]), 
	.A(sboxw[22]));
   NAND2X1 U1614 (.Y(n326), 
	.B(sboxw[7]), 
	.A(sboxw[6]));
   INVX1 U1624 (.Y(n160), 
	.A(sboxw[5]));
   INVX1 U1626 (.Y(n128), 
	.A(sboxw[29]));
endmodule

module aes_core (
	clk, 
	reset_n, 
	init, 
	next, 
	ready, 
	key, 
	block, 
	result, 
	FE_OFN37_reset_n, 
	FE_OFN38_reset_n, 
	FE_OFN39_reset_n, 
	FE_OFN40_reset_n, 
	FE_OFN42_reset_n, 
	FE_OFN43_reset_n, 
	FE_OFN44_reset_n, 
	FE_OFN45_reset_n, 
	FE_OFN46_reset_n, 
	FE_OFN47_reset_n, 
	FE_OFN48_reset_n, 
	FE_OFN49_reset_n, 
	FE_OFN50_reset_n, 
	FE_OFN51_reset_n, 
	FE_OFN53_reset_n, 
	FE_OFN54_reset_n, 
	FE_OFN55_reset_n, 
	FE_OFN56_reset_n, 
	FE_OFN58_reset_n, 
	clk_48Mhz__L6_N1, 
	clk_48Mhz__L6_N10, 
	clk_48Mhz__L6_N11, 
	clk_48Mhz__L6_N12, 
	clk_48Mhz__L6_N13, 
	clk_48Mhz__L6_N14, 
	clk_48Mhz__L6_N15, 
	clk_48Mhz__L6_N16, 
	clk_48Mhz__L6_N17, 
	clk_48Mhz__L6_N18, 
	clk_48Mhz__L6_N19, 
	clk_48Mhz__L6_N2, 
	clk_48Mhz__L6_N20, 
	clk_48Mhz__L6_N21, 
	clk_48Mhz__L6_N22, 
	clk_48Mhz__L6_N23, 
	clk_48Mhz__L6_N24, 
	clk_48Mhz__L6_N25, 
	clk_48Mhz__L6_N26, 
	clk_48Mhz__L6_N27, 
	clk_48Mhz__L6_N28, 
	clk_48Mhz__L6_N29, 
	clk_48Mhz__L6_N3, 
	clk_48Mhz__L6_N30, 
	clk_48Mhz__L6_N31, 
	clk_48Mhz__L6_N32, 
	clk_48Mhz__L6_N33, 
	clk_48Mhz__L6_N34, 
	clk_48Mhz__L6_N35, 
	clk_48Mhz__L6_N36, 
	clk_48Mhz__L6_N37, 
	clk_48Mhz__L6_N38, 
	clk_48Mhz__L6_N39, 
	clk_48Mhz__L6_N4, 
	clk_48Mhz__L6_N40, 
	clk_48Mhz__L6_N41, 
	clk_48Mhz__L6_N42, 
	clk_48Mhz__L6_N43, 
	clk_48Mhz__L6_N44, 
	clk_48Mhz__L6_N45, 
	clk_48Mhz__L6_N46, 
	clk_48Mhz__L6_N47, 
	clk_48Mhz__L6_N5, 
	clk_48Mhz__L6_N6, 
	clk_48Mhz__L6_N7, 
	clk_48Mhz__L6_N8, 
	clk_48Mhz__L6_N9);
   input clk;
   input reset_n;
   input init;
   input next;
   output ready;
   input [127:0] key;
   input [127:0] block;
   output [127:0] result;
   input FE_OFN37_reset_n;
   input FE_OFN38_reset_n;
   input FE_OFN39_reset_n;
   input FE_OFN40_reset_n;
   input FE_OFN42_reset_n;
   input FE_OFN43_reset_n;
   input FE_OFN44_reset_n;
   input FE_OFN45_reset_n;
   input FE_OFN46_reset_n;
   input FE_OFN47_reset_n;
   input FE_OFN48_reset_n;
   input FE_OFN49_reset_n;
   input FE_OFN50_reset_n;
   input FE_OFN51_reset_n;
   input FE_OFN53_reset_n;
   input FE_OFN54_reset_n;
   input FE_OFN55_reset_n;
   input FE_OFN56_reset_n;
   input FE_OFN58_reset_n;
   input clk_48Mhz__L6_N1;
   input clk_48Mhz__L6_N10;
   input clk_48Mhz__L6_N11;
   input clk_48Mhz__L6_N12;
   input clk_48Mhz__L6_N13;
   input clk_48Mhz__L6_N14;
   input clk_48Mhz__L6_N15;
   input clk_48Mhz__L6_N16;
   input clk_48Mhz__L6_N17;
   input clk_48Mhz__L6_N18;
   input clk_48Mhz__L6_N19;
   input clk_48Mhz__L6_N2;
   input clk_48Mhz__L6_N20;
   input clk_48Mhz__L6_N21;
   input clk_48Mhz__L6_N22;
   input clk_48Mhz__L6_N23;
   input clk_48Mhz__L6_N24;
   input clk_48Mhz__L6_N25;
   input clk_48Mhz__L6_N26;
   input clk_48Mhz__L6_N27;
   input clk_48Mhz__L6_N28;
   input clk_48Mhz__L6_N29;
   input clk_48Mhz__L6_N3;
   input clk_48Mhz__L6_N30;
   input clk_48Mhz__L6_N31;
   input clk_48Mhz__L6_N32;
   input clk_48Mhz__L6_N33;
   input clk_48Mhz__L6_N34;
   input clk_48Mhz__L6_N35;
   input clk_48Mhz__L6_N36;
   input clk_48Mhz__L6_N37;
   input clk_48Mhz__L6_N38;
   input clk_48Mhz__L6_N39;
   input clk_48Mhz__L6_N4;
   input clk_48Mhz__L6_N40;
   input clk_48Mhz__L6_N41;
   input clk_48Mhz__L6_N42;
   input clk_48Mhz__L6_N43;
   input clk_48Mhz__L6_N44;
   input clk_48Mhz__L6_N45;
   input clk_48Mhz__L6_N46;
   input clk_48Mhz__L6_N47;
   input clk_48Mhz__L6_N5;
   input clk_48Mhz__L6_N6;
   input clk_48Mhz__L6_N7;
   input clk_48Mhz__L6_N8;
   input clk_48Mhz__L6_N9;

   // Internal wires
   wire FE_PHN5159_n78;
   wire FE_PHN5070_ready;
   wire FE_PHN2894_n89;
   wire FE_PHN2802_ready;
   wire FE_PHN905_n78;
   wire FE_PHN820_n76;
   wire FE_PHN434_n39;
   wire FE_PHN370_n77;
   wire FE_PHN291_aes_core_ctrl_reg_1_;
   wire enc_ready;
   wire key_ready;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n84;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire [3:0] enc_round_nr;
   wire [127:0] round_key;
   wire [31:0] enc_sboxw;
   wire [31:0] new_sboxw;
   wire [31:0] keymem_sboxw;
   wire [1:0] aes_core_ctrl_reg;

   CLKBUFX1 FE_PHC5159_n78 (.Y(FE_PHN5159_n78), 
	.A(n78));
   DLY3X1 FE_PHC5070_ready (.Y(FE_PHN5070_ready), 
	.A(FE_PHN2802_ready));
   DLY3X1 FE_PHC2894_n89 (.Y(FE_PHN2894_n89), 
	.A(n89));
   DLY4X1 FE_PHC2802_ready (.Y(ready), 
	.A(FE_PHN5070_ready));
   DLY4X1 FE_PHC905_n78 (.Y(FE_PHN905_n78), 
	.A(FE_PHN5159_n78));
   DLY4X1 FE_PHC820_n76 (.Y(FE_PHN820_n76), 
	.A(n76));
   DLY4X1 FE_PHC434_n39 (.Y(FE_PHN434_n39), 
	.A(n39));
   DLY4X1 FE_PHC370_n77 (.Y(FE_PHN370_n77), 
	.A(n77));
   DLY4X1 FE_PHC291_aes_core_ctrl_reg_1_ (.Y(FE_PHN291_aes_core_ctrl_reg_1_), 
	.A(aes_core_ctrl_reg[1]));
   DFFSX1 ready_reg_reg (.SN(FE_OFN39_reset_n), 
	.QN(), 
	.Q(FE_PHN2802_ready), 
	.D(FE_PHN820_n76), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 aes_core_ctrl_reg_reg_0_ (.RN(FE_OFN39_reset_n), 
	.Q(aes_core_ctrl_reg[0]), 
	.D(FE_PHN905_n78), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 aes_core_ctrl_reg_reg_1_ (.RN(FE_OFN39_reset_n), 
	.Q(aes_core_ctrl_reg[1]), 
	.D(FE_PHN370_n77), 
	.CK(clk_48Mhz__L6_N36));
   CLKINVX3 U14 (.Y(n84), 
	.A(n44));
   INVX1 U15 (.Y(n88), 
	.A(n40));
   NAND2X1 U17 (.Y(n40), 
	.B(n90), 
	.A(FE_PHN2894_n89));
   INVX1 U18 (.Y(n87), 
	.A(n41));
   INVX1 U19 (.Y(n31), 
	.A(n55));
   AOI22X1 U20 (.Y(n55), 
	.B1(n84), 
	.B0(keymem_sboxw[28]), 
	.A1(n44), 
	.A0(enc_sboxw[28]));
   INVX1 U21 (.Y(n23), 
	.A(n63));
   AOI22X1 U22 (.Y(n63), 
	.B1(n84), 
	.B0(keymem_sboxw[20]), 
	.A1(n44), 
	.A0(enc_sboxw[20]));
   INVX1 U23 (.Y(n7), 
	.A(n49));
   AOI22X1 U24 (.Y(n49), 
	.B1(n84), 
	.B0(keymem_sboxw[4]), 
	.A1(n44), 
	.A0(enc_sboxw[4]));
   INVX1 U25 (.Y(n27), 
	.A(n59));
   AOI22X1 U26 (.Y(n59), 
	.B1(n84), 
	.B0(keymem_sboxw[24]), 
	.A1(n44), 
	.A0(enc_sboxw[24]));
   INVX1 U27 (.Y(n11), 
	.A(n45));
   AOI22X1 U28 (.Y(n45), 
	.B1(n84), 
	.B0(keymem_sboxw[8]), 
	.A1(n44), 
	.A0(enc_sboxw[8]));
   INVX1 U29 (.Y(n13), 
	.A(n74));
   AOI22X1 U30 (.Y(n74), 
	.B1(n84), 
	.B0(keymem_sboxw[10]), 
	.A1(n44), 
	.A0(enc_sboxw[10]));
   INVX1 U31 (.Y(n21), 
	.A(n66));
   AOI22X1 U32 (.Y(n66), 
	.B1(n84), 
	.B0(keymem_sboxw[18]), 
	.A1(n44), 
	.A0(enc_sboxw[18]));
   INVX1 U33 (.Y(n5), 
	.A(n53));
   AOI22X1 U34 (.Y(n53), 
	.B1(n84), 
	.B0(keymem_sboxw[2]), 
	.A1(n44), 
	.A0(enc_sboxw[2]));
   INVX1 U35 (.Y(n15), 
	.A(n72));
   AOI22X1 U36 (.Y(n72), 
	.B1(n84), 
	.B0(keymem_sboxw[12]), 
	.A1(n44), 
	.A0(enc_sboxw[12]));
   INVX1 U37 (.Y(n28), 
	.A(n58));
   AOI22X1 U38 (.Y(n58), 
	.B1(n84), 
	.B0(keymem_sboxw[25]), 
	.A1(n44), 
	.A0(enc_sboxw[25]));
   INVX1 U39 (.Y(n19), 
	.A(n68));
   AOI22X1 U40 (.Y(n68), 
	.B1(n84), 
	.B0(keymem_sboxw[16]), 
	.A1(n44), 
	.A0(enc_sboxw[16]));
   INVX1 U41 (.Y(n3), 
	.A(n75));
   AOI22X1 U42 (.Y(n75), 
	.B1(n84), 
	.B0(keymem_sboxw[0]), 
	.A1(n44), 
	.A0(enc_sboxw[0]));
   INVX1 U43 (.Y(n20), 
	.A(n67));
   AOI22X1 U44 (.Y(n67), 
	.B1(n84), 
	.B0(keymem_sboxw[17]), 
	.A1(n44), 
	.A0(enc_sboxw[17]));
   INVX1 U45 (.Y(n4), 
	.A(n64));
   AOI22X1 U46 (.Y(n64), 
	.B1(n84), 
	.B0(keymem_sboxw[1]), 
	.A1(n44), 
	.A0(enc_sboxw[1]));
   INVX1 U47 (.Y(n12), 
	.A(n43));
   AOI22X1 U48 (.Y(n43), 
	.B1(n84), 
	.B0(keymem_sboxw[9]), 
	.A1(n44), 
	.A0(enc_sboxw[9]));
   INVX1 U49 (.Y(n14), 
	.A(n73));
   AOI22X1 U50 (.Y(n73), 
	.B1(n84), 
	.B0(keymem_sboxw[11]), 
	.A1(n44), 
	.A0(enc_sboxw[11]));
   INVX1 U51 (.Y(n30), 
	.A(n56));
   AOI22X1 U52 (.Y(n56), 
	.B1(n84), 
	.B0(keymem_sboxw[27]), 
	.A1(n44), 
	.A0(enc_sboxw[27]));
   INVX1 U53 (.Y(n22), 
	.A(n65));
   AOI22X1 U54 (.Y(n65), 
	.B1(n84), 
	.B0(keymem_sboxw[19]), 
	.A1(n44), 
	.A0(enc_sboxw[19]));
   INVX1 U55 (.Y(n6), 
	.A(n50));
   AOI22X1 U56 (.Y(n50), 
	.B1(n84), 
	.B0(keymem_sboxw[3]), 
	.A1(n44), 
	.A0(enc_sboxw[3]));
   INVX1 U57 (.Y(n8), 
	.A(n48));
   AOI22X1 U58 (.Y(n48), 
	.B1(n84), 
	.B0(keymem_sboxw[5]), 
	.A1(n44), 
	.A0(enc_sboxw[5]));
   AOI22X1 U60 (.Y(n71), 
	.B1(n84), 
	.B0(keymem_sboxw[13]), 
	.A1(n44), 
	.A0(enc_sboxw[13]));
   INVX1 U61 (.Y(n32), 
	.A(n54));
   AOI22X1 U62 (.Y(n54), 
	.B1(n84), 
	.B0(keymem_sboxw[29]), 
	.A1(n44), 
	.A0(enc_sboxw[29]));
   INVX1 U63 (.Y(n24), 
	.A(n62));
   AOI22X1 U64 (.Y(n62), 
	.B1(n84), 
	.B0(keymem_sboxw[21]), 
	.A1(n44), 
	.A0(enc_sboxw[21]));
   OAI21X2 U65 (.Y(n44), 
	.B0(n90), 
	.A1(init), 
	.A0(aes_core_ctrl_reg[0]));
   INVX1 U66 (.Y(n90), 
	.A(FE_PHN291_aes_core_ctrl_reg_1_));
   INVX1 U67 (.Y(n29), 
	.A(n57));
   AOI22X1 U68 (.Y(n57), 
	.B1(n84), 
	.B0(keymem_sboxw[26]), 
	.A1(n44), 
	.A0(enc_sboxw[26]));
   INVX1 U69 (.Y(n25), 
	.A(n61));
   AOI22X1 U70 (.Y(n61), 
	.B1(n84), 
	.B0(keymem_sboxw[22]), 
	.A1(n44), 
	.A0(enc_sboxw[22]));
   INVX1 U71 (.Y(n9), 
	.A(n47));
   AOI22X1 U72 (.Y(n47), 
	.B1(n84), 
	.B0(keymem_sboxw[6]), 
	.A1(n44), 
	.A0(enc_sboxw[6]));
   INVX1 U73 (.Y(n33), 
	.A(n52));
   AOI22X1 U74 (.Y(n52), 
	.B1(n84), 
	.B0(keymem_sboxw[30]), 
	.A1(n44), 
	.A0(enc_sboxw[30]));
   INVX1 U75 (.Y(n17), 
	.A(n70));
   AOI22X1 U76 (.Y(n70), 
	.B1(n84), 
	.B0(keymem_sboxw[14]), 
	.A1(n44), 
	.A0(enc_sboxw[14]));
   INVX1 U77 (.Y(n18), 
	.A(n69));
   AOI22X1 U78 (.Y(n69), 
	.B1(n84), 
	.B0(keymem_sboxw[15]), 
	.A1(n44), 
	.A0(enc_sboxw[15]));
   INVX1 U79 (.Y(n26), 
	.A(n60));
   AOI22X1 U80 (.Y(n60), 
	.B1(n84), 
	.B0(keymem_sboxw[23]), 
	.A1(n44), 
	.A0(enc_sboxw[23]));
   INVX1 U81 (.Y(n34), 
	.A(n51));
   AOI22X1 U82 (.Y(n51), 
	.B1(n84), 
	.B0(keymem_sboxw[31]), 
	.A1(n44), 
	.A0(enc_sboxw[31]));
   INVX1 U83 (.Y(n10), 
	.A(n46));
   AOI22X1 U84 (.Y(n46), 
	.B1(n84), 
	.B0(keymem_sboxw[7]), 
	.A1(n44), 
	.A0(enc_sboxw[7]));
   AOI33X1 U85 (.Y(n39), 
	.B2(key_ready), 
	.B1(n90), 
	.B0(aes_core_ctrl_reg[0]), 
	.A2(enc_ready), 
	.A1(n89), 
	.A0(FE_PHN291_aes_core_ctrl_reg_1_));
   OAI32X1 U86 (.Y(n77), 
	.B1(n41), 
	.B0(n90), 
	.A2(n87), 
	.A1(init), 
	.A0(n40));
   INVX1 U87 (.Y(n89), 
	.A(aes_core_ctrl_reg[0]));
   NAND2X1 U88 (.Y(n41), 
	.B(n42), 
	.A(FE_PHN434_n39));
   OAI21XL U89 (.Y(n42), 
	.B0(n88), 
	.A1(next), 
	.A0(init));
   OAI2BB2X1 U90 (.Y(n78), 
	.B1(n41), 
	.B0(FE_PHN2894_n89), 
	.A1N(init), 
	.A0N(n88));
   OAI2BB1X1 U91 (.Y(n76), 
	.B0(FE_PHN434_n39), 
	.A1N(n87), 
	.A0N(ready));
   aes_encipher_block enc_block (.clk(clk_48Mhz__L6_N21), 
	.reset_n(FE_OFN38_reset_n), 
	.next(next), 
	.round(enc_round_nr), 
	.round_key(round_key), 
	.sboxw(enc_sboxw), 
	.new_sboxw(new_sboxw), 
	.block(block), 
	.new_block(result), 
	.ready(enc_ready), 
	.FE_OFN39_reset_n(FE_OFN39_reset_n), 
	.FE_OFN43_reset_n(FE_OFN43_reset_n), 
	.FE_OFN49_reset_n(FE_OFN49_reset_n), 
	.FE_OFN50_reset_n(FE_OFN50_reset_n), 
	.FE_OFN51_reset_n(FE_OFN51_reset_n), 
	.FE_OFN54_reset_n(FE_OFN54_reset_n), 
	.FE_OFN55_reset_n(FE_OFN55_reset_n), 
	.FE_OFN56_reset_n(FE_OFN56_reset_n), 
	.clk_48Mhz__L6_N23(clk_48Mhz__L6_N23), 
	.clk_48Mhz__L6_N37(clk_48Mhz__L6_N37), 
	.clk_48Mhz__L6_N39(clk_48Mhz__L6_N39), 
	.clk_48Mhz__L6_N40(clk_48Mhz__L6_N40), 
	.clk_48Mhz__L6_N41(clk_48Mhz__L6_N41), 
	.clk_48Mhz__L6_N44(clk_48Mhz__L6_N44), 
	.clk_48Mhz__L6_N46(clk_48Mhz__L6_N46), 
	.clk_48Mhz__L6_N47(clk_48Mhz__L6_N47), 
	.clk_48Mhz__L6_N5(clk_48Mhz__L6_N5), 
	.clk_48Mhz__L6_N8(clk_48Mhz__L6_N8), 
	.clk_48Mhz__L6_N9(clk_48Mhz__L6_N9));
   aes_key_mem keymem (.clk(clk), 
	.reset_n(reset_n), 
	.key(key), 
	.init(init), 
	.round(enc_round_nr), 
	.round_key(round_key), 
	.ready(key_ready), 
	.sboxw(keymem_sboxw), 
	.new_sboxw(new_sboxw), 
	.FE_OFN37_reset_n(FE_OFN37_reset_n), 
	.FE_OFN39_reset_n(FE_OFN39_reset_n), 
	.FE_OFN40_reset_n(FE_OFN40_reset_n), 
	.FE_OFN42_reset_n(FE_OFN42_reset_n), 
	.FE_OFN43_reset_n(FE_OFN43_reset_n), 
	.FE_OFN44_reset_n(FE_OFN44_reset_n), 
	.FE_OFN45_reset_n(FE_OFN45_reset_n), 
	.FE_OFN46_reset_n(FE_OFN46_reset_n), 
	.FE_OFN47_reset_n(FE_OFN47_reset_n), 
	.FE_OFN48_reset_n(FE_OFN48_reset_n), 
	.FE_OFN53_reset_n(FE_OFN53_reset_n), 
	.FE_OFN55_reset_n(FE_OFN55_reset_n), 
	.FE_OFN58_reset_n(FE_OFN58_reset_n), 
	.clk_48Mhz__L6_N1(clk_48Mhz__L6_N1), 
	.clk_48Mhz__L6_N10(clk_48Mhz__L6_N10), 
	.clk_48Mhz__L6_N11(clk_48Mhz__L6_N11), 
	.clk_48Mhz__L6_N12(clk_48Mhz__L6_N12), 
	.clk_48Mhz__L6_N13(clk_48Mhz__L6_N13), 
	.clk_48Mhz__L6_N14(clk_48Mhz__L6_N14), 
	.clk_48Mhz__L6_N15(clk_48Mhz__L6_N15), 
	.clk_48Mhz__L6_N16(clk_48Mhz__L6_N16), 
	.clk_48Mhz__L6_N17(clk_48Mhz__L6_N17), 
	.clk_48Mhz__L6_N18(clk_48Mhz__L6_N18), 
	.clk_48Mhz__L6_N19(clk_48Mhz__L6_N19), 
	.clk_48Mhz__L6_N2(clk_48Mhz__L6_N2), 
	.clk_48Mhz__L6_N20(clk_48Mhz__L6_N20), 
	.clk_48Mhz__L6_N21(clk_48Mhz__L6_N21), 
	.clk_48Mhz__L6_N22(clk_48Mhz__L6_N22), 
	.clk_48Mhz__L6_N23(clk_48Mhz__L6_N23), 
	.clk_48Mhz__L6_N24(clk_48Mhz__L6_N24), 
	.clk_48Mhz__L6_N25(clk_48Mhz__L6_N25), 
	.clk_48Mhz__L6_N26(clk_48Mhz__L6_N26), 
	.clk_48Mhz__L6_N27(clk_48Mhz__L6_N27), 
	.clk_48Mhz__L6_N28(clk_48Mhz__L6_N28), 
	.clk_48Mhz__L6_N29(clk_48Mhz__L6_N29), 
	.clk_48Mhz__L6_N3(clk_48Mhz__L6_N3), 
	.clk_48Mhz__L6_N30(clk_48Mhz__L6_N30), 
	.clk_48Mhz__L6_N31(clk_48Mhz__L6_N31), 
	.clk_48Mhz__L6_N32(clk_48Mhz__L6_N32), 
	.clk_48Mhz__L6_N33(clk_48Mhz__L6_N33), 
	.clk_48Mhz__L6_N34(clk_48Mhz__L6_N34), 
	.clk_48Mhz__L6_N35(clk_48Mhz__L6_N35), 
	.clk_48Mhz__L6_N36(clk_48Mhz__L6_N36), 
	.clk_48Mhz__L6_N37(clk_48Mhz__L6_N37), 
	.clk_48Mhz__L6_N38(clk_48Mhz__L6_N38), 
	.clk_48Mhz__L6_N4(clk_48Mhz__L6_N4), 
	.clk_48Mhz__L6_N42(clk_48Mhz__L6_N42), 
	.clk_48Mhz__L6_N43(clk_48Mhz__L6_N43), 
	.clk_48Mhz__L6_N44(clk_48Mhz__L6_N44), 
	.clk_48Mhz__L6_N45(clk_48Mhz__L6_N45), 
	.clk_48Mhz__L6_N46(clk_48Mhz__L6_N46), 
	.clk_48Mhz__L6_N47(clk_48Mhz__L6_N47), 
	.clk_48Mhz__L6_N5(clk_48Mhz__L6_N5), 
	.clk_48Mhz__L6_N6(clk_48Mhz__L6_N6), 
	.clk_48Mhz__L6_N7(clk_48Mhz__L6_N7), 
	.clk_48Mhz__L6_N8(clk_48Mhz__L6_N8), 
	.clk_48Mhz__L6_N9(clk_48Mhz__L6_N9));
   aes_sbox sbox_inst (.sboxw({ n34,
		n33,
		n32,
		n31,
		n30,
		n29,
		n28,
		n27,
		n26,
		n25,
		n24,
		n23,
		n22,
		n21,
		n20,
		n19,
		n18,
		n17,
		n71,
		n15,
		n14,
		n13,
		n12,
		n11,
		n10,
		n9,
		n8,
		n7,
		n6,
		n5,
		n4,
		n3 }), 
	.new_sboxw(new_sboxw));
endmodule

module reg_in (
	reset_n, 
	clk_48Mhz, 
	plain_byte_in, 
	plain_byte_valid, 
	plain_finish, 
	plain_key_out, 
	FE_OFN38_reset_n, 
	FE_OFN39_reset_n, 
	FE_OFN40_reset_n, 
	FE_OFN42_reset_n, 
	FE_OFN43_reset_n, 
	FE_OFN44_reset_n, 
	FE_OFN45_reset_n, 
	FE_OFN47_reset_n, 
	FE_OFN49_reset_n, 
	FE_OFN50_reset_n, 
	FE_OFN51_reset_n, 
	FE_OFN55_reset_n, 
	FE_OFN56_reset_n, 
	FE_OFN58_reset_n, 
	clk_48Mhz__L6_N1, 
	clk_48Mhz__L6_N10, 
	clk_48Mhz__L6_N11, 
	clk_48Mhz__L6_N14, 
	clk_48Mhz__L6_N15, 
	clk_48Mhz__L6_N2, 
	clk_48Mhz__L6_N20, 
	clk_48Mhz__L6_N21, 
	clk_48Mhz__L6_N23, 
	clk_48Mhz__L6_N25, 
	clk_48Mhz__L6_N27, 
	clk_48Mhz__L6_N28, 
	clk_48Mhz__L6_N29, 
	clk_48Mhz__L6_N35, 
	clk_48Mhz__L6_N37, 
	clk_48Mhz__L6_N39, 
	clk_48Mhz__L6_N4, 
	clk_48Mhz__L6_N40, 
	clk_48Mhz__L6_N41, 
	clk_48Mhz__L6_N5, 
	clk_48Mhz__L6_N6, 
	clk_48Mhz__L6_N8, 
	clk_48Mhz__L6_N9);
   input reset_n;
   input clk_48Mhz;
   input [7:0] plain_byte_in;
   input plain_byte_valid;
   input plain_finish;
   output [255:0] plain_key_out;
   input FE_OFN38_reset_n;
   input FE_OFN39_reset_n;
   input FE_OFN40_reset_n;
   input FE_OFN42_reset_n;
   input FE_OFN43_reset_n;
   input FE_OFN44_reset_n;
   input FE_OFN45_reset_n;
   input FE_OFN47_reset_n;
   input FE_OFN49_reset_n;
   input FE_OFN50_reset_n;
   input FE_OFN51_reset_n;
   input FE_OFN55_reset_n;
   input FE_OFN56_reset_n;
   input FE_OFN58_reset_n;
   input clk_48Mhz__L6_N1;
   input clk_48Mhz__L6_N10;
   input clk_48Mhz__L6_N11;
   input clk_48Mhz__L6_N14;
   input clk_48Mhz__L6_N15;
   input clk_48Mhz__L6_N2;
   input clk_48Mhz__L6_N20;
   input clk_48Mhz__L6_N21;
   input clk_48Mhz__L6_N23;
   input clk_48Mhz__L6_N25;
   input clk_48Mhz__L6_N27;
   input clk_48Mhz__L6_N28;
   input clk_48Mhz__L6_N29;
   input clk_48Mhz__L6_N35;
   input clk_48Mhz__L6_N37;
   input clk_48Mhz__L6_N39;
   input clk_48Mhz__L6_N4;
   input clk_48Mhz__L6_N40;
   input clk_48Mhz__L6_N41;
   input clk_48Mhz__L6_N5;
   input clk_48Mhz__L6_N6;
   input clk_48Mhz__L6_N8;
   input clk_48Mhz__L6_N9;

   // Internal wires
   wire FE_PHN5257_plain_text_28_;
   wire FE_PHN5255_plain_text_185_;
   wire FE_PHN5254_n505;
   wire FE_PHN5243_plain_text_78_;
   wire FE_PHN5242_plain_text_12_;
   wire FE_PHN5241_n505;
   wire FE_PHN5240_plain_text_185_;
   wire FE_PHN5239_plain_text_153_;
   wire FE_PHN5238_n484;
   wire FE_PHN5237_n420;
   wire FE_PHN5236_plain_text_106_;
   wire FE_PHN5234_plain_text_121_;
   wire FE_PHN5232_n516;
   wire FE_PHN5231_plain_text_49_;
   wire FE_PHN5230_Din_241_;
   wire FE_PHN5171_plain_text_49_;
   wire FE_PHN5170_plain_text_1_;
   wire FE_PHN5158_n502;
   wire FE_PHN5157_n516;
   wire FE_PHN5156_plain_text_49_;
   wire FE_PHN5155_plain_text_1_;
   wire FE_PHN5154_plain_text_121_;
   wire FE_PHN5072_plain_text_125_;
   wire FE_PHN5069_pf0;
   wire FE_PHN5067_pbv0;
   wire FE_PHN5048_n475;
   wire FE_PHN5046_n474;
   wire FE_PHN3610_n265;
   wire FE_PHN3609_n383;
   wire FE_PHN3608_n262;
   wire FE_PHN3607_plain_text_235_;
   wire FE_PHN3606_n261;
   wire FE_PHN3605_n285;
   wire FE_PHN3604_n399;
   wire FE_PHN3603_n442;
   wire FE_PHN3602_n417;
   wire FE_PHN3601_n382;
   wire FE_PHN3600_n407;
   wire FE_PHN3599_n329;
   wire FE_PHN3598_n470;
   wire FE_PHN3597_plain_text_172_;
   wire FE_PHN3596_n270;
   wire FE_PHN3595_n278;
   wire FE_PHN3594_n284;
   wire FE_PHN3593_n271;
   wire FE_PHN3592_n267;
   wire FE_PHN3591_n277;
   wire FE_PHN3590_n409;
   wire FE_PHN3589_n260;
   wire FE_PHN3588_plain_text_204_;
   wire FE_PHN3587_n319;
   wire FE_PHN3586_n264;
   wire FE_PHN3585_n318;
   wire FE_PHN3584_n263;
   wire FE_PHN3583_n314;
   wire FE_PHN3582_n488;
   wire FE_PHN3581_n351;
   wire FE_PHN3580_n506;
   wire FE_PHN3579_n367;
   wire FE_PHN3578_n266;
   wire FE_PHN3577_n288;
   wire FE_PHN3576_plain_text_139_;
   wire FE_PHN3575_n378;
   wire FE_PHN3574_n472;
   wire FE_PHN3573_n372;
   wire FE_PHN3572_n374;
   wire FE_PHN3571_n448;
   wire FE_PHN3570_n415;
   wire FE_PHN3569_n381;
   wire FE_PHN3568_n449;
   wire FE_PHN3567_n295;
   wire FE_PHN3566_n331;
   wire FE_PHN3565_n316;
   wire FE_PHN3564_n333;
   wire FE_PHN3563_n353;
   wire FE_PHN3562_n274;
   wire FE_PHN3561_n462;
   wire FE_PHN3560_n380;
   wire FE_PHN3559_plain_text_12_;
   wire FE_PHN3558_n439;
   wire FE_PHN3557_n328;
   wire FE_PHN3556_n317;
   wire FE_PHN3555_n406;
   wire FE_PHN3554_n468;
   wire FE_PHN3553_n369;
   wire FE_PHN3552_n273;
   wire FE_PHN3551_n289;
   wire FE_PHN3550_n401;
   wire FE_PHN3549_n416;
   wire FE_PHN3548_n339;
   wire FE_PHN3547_n363;
   wire FE_PHN3546_n345;
   wire FE_PHN3545_n460;
   wire FE_PHN3544_n446;
   wire FE_PHN3543_n300;
   wire FE_PHN3542_n355;
   wire FE_PHN3541_n365;
   wire FE_PHN3540_n361;
   wire FE_PHN3539_n438;
   wire FE_PHN3538_n349;
   wire FE_PHN3537_n390;
   wire FE_PHN3536_n292;
   wire FE_PHN3535_n275;
   wire FE_PHN3534_n463;
   wire FE_PHN3533_n330;
   wire FE_PHN3532_n337;
   wire FE_PHN3531_n375;
   wire FE_PHN3530_n282;
   wire FE_PHN3529_n394;
   wire FE_PHN3528_n308;
   wire FE_PHN3527_n326;
   wire FE_PHN3526_n366;
   wire FE_PHN3525_n344;
   wire FE_PHN3524_n352;
   wire FE_PHN3523_n362;
   wire FE_PHN3522_n307;
   wire FE_PHN3521_n342;
   wire FE_PHN3520_n303;
   wire FE_PHN3519_n348;
   wire FE_PHN3518_n485;
   wire FE_PHN3517_n503;
   wire FE_PHN3516_n371;
   wire FE_PHN3515_n296;
   wire FE_PHN3514_n477;
   wire FE_PHN3513_n405;
   wire FE_PHN3512_n334;
   wire FE_PHN3511_n433;
   wire FE_PHN3510_n357;
   wire FE_PHN3509_n321;
   wire FE_PHN3508_n441;
   wire FE_PHN3507_n276;
   wire FE_PHN3506_n400;
   wire FE_PHN3505_n341;
   wire FE_PHN3504_n496;
   wire FE_PHN3503_n354;
   wire FE_PHN3502_n280;
   wire FE_PHN3501_n324;
   wire FE_PHN3500_n379;
   wire FE_PHN3499_n454;
   wire FE_PHN3498_n482;
   wire FE_PHN3497_n480;
   wire FE_PHN3496_n325;
   wire FE_PHN3495_n450;
   wire FE_PHN3494_n473;
   wire FE_PHN3493_n452;
   wire FE_PHN3492_n440;
   wire FE_PHN3491_n320;
   wire FE_PHN3490_n279;
   wire FE_PHN3489_n286;
   wire FE_PHN3488_n297;
   wire FE_PHN3487_n364;
   wire FE_PHN3486_n350;
   wire FE_PHN3485_n310;
   wire FE_PHN3484_n347;
   wire FE_PHN3483_n359;
   wire FE_PHN3482_n312;
   wire FE_PHN3481_n304;
   wire FE_PHN3480_n302;
   wire FE_PHN3479_n343;
   wire FE_PHN3478_n465;
   wire FE_PHN3477_n311;
   wire FE_PHN3476_n346;
   wire FE_PHN3475_n293;
   wire FE_PHN3474_n306;
   wire FE_PHN3473_n338;
   wire FE_PHN3472_n373;
   wire FE_PHN3471_n428;
   wire FE_PHN3470_n499;
   wire FE_PHN3469_n269;
   wire FE_PHN3468_n429;
   wire FE_PHN3467_n309;
   wire FE_PHN3466_n393;
   wire FE_PHN3465_n340;
   wire FE_PHN3464_n268;
   wire FE_PHN3463_n305;
   wire FE_PHN3462_n476;
   wire FE_PHN3461_n335;
   wire FE_PHN3460_n421;
   wire FE_PHN3459_n368;
   wire FE_PHN3458_n356;
   wire FE_PHN3457_n389;
   wire FE_PHN3456_n332;
   wire FE_PHN3455_n453;
   wire FE_PHN3454_n392;
   wire FE_PHN3453_n322;
   wire FE_PHN3452_n294;
   wire FE_PHN3451_n391;
   wire FE_PHN3450_n336;
   wire FE_PHN3449_n358;
   wire FE_PHN3448_n388;
   wire FE_PHN3447_n403;
   wire FE_PHN3446_n360;
   wire FE_PHN3445_n500;
   wire FE_PHN3443_n483;
   wire FE_PHN3442_n398;
   wire FE_PHN3441_n431;
   wire FE_PHN3440_n430;
   wire FE_PHN3439_n461;
   wire FE_PHN3438_n299;
   wire FE_PHN3436_n397;
   wire FE_PHN3432_n313;
   wire FE_PHN3405_n491;
   wire FE_PHN3404_plain_text_32_;
   wire FE_PHN3402_n410;
   wire FE_PHN3401_n419;
   wire FE_PHN3400_plain_text_42_;
   wire FE_PHN3399_n418;
   wire FE_PHN3398_n323;
   wire FE_PHN3397_n467;
   wire FE_PHN3396_n411;
   wire FE_PHN3395_n466;
   wire FE_PHN3394_n490;
   wire FE_PHN3393_n435;
   wire FE_PHN3392_n458;
   wire FE_PHN3391_plain_text_0_;
   wire FE_PHN3390_plain_text_147_;
   wire FE_PHN3389_plain_text_157_;
   wire FE_PHN3387_n624;
   wire FE_PHN3386_plain_text_133_;
   wire FE_PHN3385_n620;
   wire FE_PHN3384_n709;
   wire FE_PHN3383_n724;
   wire FE_PHN3382_plain_text_18_;
   wire FE_PHN3381_n686;
   wire FE_PHN3380_n638;
   wire FE_PHN3379_plain_text_33_;
   wire FE_PHN3377_n542;
   wire FE_PHN3376_plain_text_59_;
   wire FE_PHN3375_n545;
   wire FE_PHN3374_n584;
   wire FE_PHN3372_n543;
   wire FE_PHN3370_n658;
   wire FE_PHN3369_plain_text_146_;
   wire FE_PHN3368_n608;
   wire FE_PHN3367_plain_text_196_;
   wire FE_PHN3366_n605;
   wire FE_PHN3364_n582;
   wire FE_PHN3363_plain_text_163_;
   wire FE_PHN3361_n693;
   wire FE_PHN3357_n519;
   wire FE_PHN3355_plain_text_225_;
   wire FE_PHN3354_plain_text_168_;
   wire FE_PHN3352_n617;
   wire FE_PHN3350_plain_text_203_;
   wire FE_PHN3348_plain_text_52_;
   wire FE_PHN3347_n736;
   wire FE_PHN3346_n557;
   wire FE_PHN3337_plain_text_241_;
   wire FE_PHN3336_plain_text_243_;
   wire FE_PHN3320_plain_text_55_;
   wire FE_PHN3318_plain_text_23_;
   wire FE_PHN3317_n768;
   wire FE_PHN3311_plain_text_193_;
   wire FE_PHN3306_n726;
   wire FE_PHN3300_n612;
   wire FE_PHN3299_plain_text_31_;
   wire FE_PHN3298_plain_text_161_;
   wire FE_PHN3297_n558;
   wire FE_PHN3291_n741;
   wire FE_PHN3287_plain_text_192_;
   wire FE_PHN3286_n522;
   wire FE_PHN3280_plain_text_21_;
   wire FE_PHN3279_n704;
   wire FE_PHN3264_n645;
   wire FE_PHN3257_n661;
   wire FE_PHN3254_n765;
   wire FE_PHN3199_n606;
   wire FE_PHN3182_plain_text_1_;
   wire FE_PHN3181_plain_text_2_;
   wire FE_PHN3176_plain_text_123_;
   wire FE_PHN3175_plain_text_6_;
   wire FE_PHN3174_plain_text_14_;
   wire FE_PHN3172_n717;
   wire FE_PHN3171_plain_text_7_;
   wire FE_PHN3170_n771;
   wire FE_PHN3169_plain_text_182_;
   wire FE_PHN3168_n716;
   wire FE_PHN3167_plain_text_122_;
   wire FE_PHN3166_plain_text_179_;
   wire FE_PHN3165_plain_text_25_;
   wire FE_PHN3164_plain_text_69_;
   wire FE_PHN3163_plain_text_11_;
   wire FE_PHN3162_plain_text_228_;
   wire FE_PHN3159_n744;
   wire FE_PHN3158_n712;
   wire FE_PHN3157_plain_text_231_;
   wire FE_PHN3156_plain_text_171_;
   wire FE_PHN3155_n723;
   wire FE_PHN3154_plain_text_189_;
   wire FE_PHN3153_plain_text_205_;
   wire FE_PHN3152_plain_text_210_;
   wire FE_PHN3151_plain_text_48_;
   wire FE_PHN3150_n746;
   wire FE_PHN3148_plain_text_178_;
   wire FE_PHN3147_plain_text_28_;
   wire FE_PHN3146_plain_text_65_;
   wire FE_PHN3145_n748;
   wire FE_PHN3144_n713;
   wire FE_PHN3143_plain_text_206_;
   wire FE_PHN3142_n641;
   wire FE_PHN3141_plain_text_54_;
   wire FE_PHN3140_n714;
   wire FE_PHN3139_plain_text_198_;
   wire FE_PHN3138_n715;
   wire FE_PHN3137_plain_text_138_;
   wire FE_PHN3136_plain_text_216_;
   wire FE_PHN3135_plain_text_56_;
   wire FE_PHN3134_n525;
   wire FE_PHN3133_plain_text_170_;
   wire FE_PHN3132_n539;
   wire FE_PHN3131_plain_text_169_;
   wire FE_PHN3130_n745;
   wire FE_PHN3129_n750;
   wire FE_PHN3128_plain_text_81_;
   wire FE_PHN3127_n754;
   wire FE_PHN3126_plain_text_141_;
   wire FE_PHN3125_plain_text_68_;
   wire FE_PHN3124_plain_text_72_;
   wire FE_PHN3123_n537;
   wire FE_PHN3122_n530;
   wire FE_PHN3121_plain_text_128_;
   wire FE_PHN3120_n751;
   wire FE_PHN3119_n743;
   wire FE_PHN3118_n722;
   wire FE_PHN3117_n749;
   wire FE_PHN3116_plain_text_175_;
   wire FE_PHN3115_n719;
   wire FE_PHN3114_plain_text_137_;
   wire FE_PHN3113_n562;
   wire FE_PHN3112_plain_text_129_;
   wire FE_PHN3111_n640;
   wire FE_PHN3110_plain_text_47_;
   wire FE_PHN3109_n538;
   wire FE_PHN3103_plain_text_10_;
   wire FE_PHN3102_plain_text_118_;
   wire FE_PHN3101_plain_text_227_;
   wire FE_PHN3100_plain_text_212_;
   wire FE_PHN3099_plain_text_162_;
   wire FE_PHN3098_plain_text_60_;
   wire FE_PHN3097_plain_text_150_;
   wire FE_PHN3096_plain_text_234_;
   wire FE_PHN3093_plain_text_217_;
   wire FE_PHN3092_plain_text_75_;
   wire FE_PHN3090_plain_text_49_;
   wire FE_PHN3088_plain_text_251_;
   wire FE_PHN3087_plain_text_254_;
   wire FE_PHN3086_plain_text_180_;
   wire FE_PHN3084_plain_text_191_;
   wire FE_PHN3083_plain_text_46_;
   wire FE_PHN3082_plain_text_249_;
   wire FE_PHN3080_n384;
   wire FE_PHN3079_plain_text_5_;
   wire FE_PHN3078_n479;
   wire FE_PHN3077_n414;
   wire FE_PHN3076_n447;
   wire FE_PHN3075_n298;
   wire FE_PHN3074_plain_text_3_;
   wire FE_PHN3073_n420;
   wire FE_PHN3072_n437;
   wire FE_PHN3071_n478;
   wire FE_PHN3070_n481;
   wire FE_PHN3069_n445;
   wire FE_PHN3068_n413;
   wire FE_PHN3067_n376;
   wire FE_PHN3066_n301;
   wire FE_PHN3065_plain_text_246_;
   wire FE_PHN3064_n377;
   wire FE_PHN3063_plain_text_58_;
   wire FE_PHN3062_n412;
   wire FE_PHN3061_n327;
   wire FE_PHN3060_n464;
   wire FE_PHN3059_n455;
   wire FE_PHN3058_n436;
   wire FE_PHN3057_n290;
   wire FE_PHN3056_n487;
   wire FE_PHN3055_n504;
   wire FE_PHN3054_plain_text_24_;
   wire FE_PHN3053_n444;
   wire FE_PHN3052_plain_text_114_;
   wire FE_PHN3051_plain_text_93_;
   wire FE_PHN3050_n515;
   wire FE_PHN3049_n497;
   wire FE_PHN3048_plain_text_73_;
   wire FE_PHN3047_n493;
   wire FE_PHN3046_n484;
   wire FE_PHN3045_plain_text_190_;
   wire FE_PHN3044_plain_text_17_;
   wire FE_PHN3043_plain_text_109_;
   wire FE_PHN3042_n287;
   wire FE_PHN3041_plain_text_95_;
   wire FE_PHN3040_plain_text_200_;
   wire FE_PHN3039_n370;
   wire FE_PHN3038_plain_text_101_;
   wire FE_PHN3037_plain_text_107_;
   wire FE_PHN3036_n489;
   wire FE_PHN3035_n471;
   wire FE_PHN3034_plain_text_29_;
   wire FE_PHN3033_plain_text_103_;
   wire FE_PHN3032_plain_text_120_;
   wire FE_PHN3031_plain_text_202_;
   wire FE_PHN3030_plain_text_112_;
   wire FE_PHN3029_plain_text_22_;
   wire FE_PHN3028_n422;
   wire FE_PHN3027_plain_text_79_;
   wire FE_PHN3026_n505;
   wire FE_PHN3025_plain_text_131_;
   wire FE_PHN3024_n502;
   wire FE_PHN3023_plain_text_207_;
   wire FE_PHN3022_n402;
   wire FE_PHN3021_n396;
   wire FE_PHN3020_plain_text_99_;
   wire FE_PHN3019_plain_text_115_;
   wire FE_PHN3018_n501;
   wire FE_PHN3017_plain_text_90_;
   wire FE_PHN3016_plain_text_121_;
   wire FE_PHN3015_plain_text_91_;
   wire FE_PHN3014_n494;
   wire FE_PHN3013_plain_text_70_;
   wire FE_PHN3012_plain_text_194_;
   wire FE_PHN3011_plain_text_61_;
   wire FE_PHN3010_plain_text_149_;
   wire FE_PHN3009_plain_text_89_;
   wire FE_PHN3008_plain_text_208_;
   wire FE_PHN3007_plain_text_156_;
   wire FE_PHN3006_plain_text_84_;
   wire FE_PHN3005_plain_text_66_;
   wire FE_PHN3004_plain_text_223_;
   wire FE_PHN3003_plain_text_159_;
   wire FE_PHN3002_plain_text_71_;
   wire FE_PHN3001_plain_text_82_;
   wire FE_PHN3000_plain_text_78_;
   wire FE_PHN2999_plain_text_57_;
   wire FE_PHN2998_plain_text_92_;
   wire FE_PHN2997_n495;
   wire FE_PHN2996_n492;
   wire FE_PHN2995_plain_text_85_;
   wire FE_PHN2994_plain_text_186_;
   wire FE_PHN2992_plain_text_98_;
   wire FE_PHN2991_plain_text_106_;
   wire FE_PHN2989_plain_text_181_;
   wire FE_PHN2988_plain_text_173_;
   wire FE_PHN2987_plain_text_86_;
   wire FE_PHN2986_n507;
   wire FE_PHN2985_plain_text_74_;
   wire FE_PHN2984_plain_text_158_;
   wire FE_PHN2981_plain_text_102_;
   wire FE_PHN2980_plain_text_94_;
   wire FE_PHN2979_plain_text_104_;
   wire FE_PHN2978_plain_text_37_;
   wire FE_PHN2977_plain_text_80_;
   wire FE_PHN2976_plain_text_164_;
   wire FE_PHN2975_n424;
   wire FE_PHN2974_n404;
   wire FE_PHN2973_plain_text_96_;
   wire FE_PHN2972_plain_text_87_;
   wire FE_PHN2971_plain_text_9_;
   wire FE_PHN2969_plain_text_213_;
   wire FE_PHN2968_plain_text_220_;
   wire FE_PHN2967_n432;
   wire FE_PHN2966_plain_text_222_;
   wire FE_PHN2965_plain_text_83_;
   wire FE_PHN2964_plain_text_148_;
   wire FE_PHN2963_n408;
   wire FE_PHN2962_n469;
   wire FE_PHN2961_plain_text_45_;
   wire FE_PHN2960_plain_text_111_;
   wire FE_PHN2959_plain_text_63_;
   wire FE_PHN2958_plain_text_88_;
   wire FE_PHN2957_plain_text_105_;
   wire FE_PHN2953_plain_text_236_;
   wire FE_PHN2952_plain_text_97_;
   wire FE_PHN2950_plain_text_44_;
   wire FE_PHN2949_plain_text_108_;
   wire FE_PHN2948_plain_text_119_;
   wire FE_PHN2945_plain_text_113_;
   wire FE_PHN2944_plain_text_76_;
   wire FE_PHN2943_plain_text_151_;
   wire FE_PHN2942_plain_text_100_;
   wire FE_PHN2940_n510;
   wire FE_PHN2939_n511;
   wire FE_PHN2938_n514;
   wire FE_PHN2937_n512;
   wire FE_PHN2934_n513;
   wire FE_PHN2933_plain_text_188_;
   wire FE_PHN2932_plain_text_34_;
   wire FE_PHN2931_n451;
   wire FE_PHN2929_plain_text_51_;
   wire FE_PHN2928_n457;
   wire FE_PHN2926_plain_text_53_;
   wire FE_PHN2925_plain_text_39_;
   wire FE_PHN2924_n509;
   wire FE_PHN2923_Din_12_;
   wire FE_PHN2922_Din_21_;
   wire FE_PHN2921_Din_23_;
   wire FE_PHN2920_Din_55_;
   wire FE_PHN2889_n575;
   wire FE_PHN2888_plain_text_4_;
   wire FE_PHN2887_plain_text_155_;
   wire FE_PHN2886_n593;
   wire FE_PHN2885_plain_text_15_;
   wire FE_PHN2884_plain_text_40_;
   wire FE_PHN2883_n626;
   wire FE_PHN2882_plain_text_77_;
   wire FE_PHN2881_n688;
   wire FE_PHN2880_plain_text_16_;
   wire FE_PHN2879_n516;
   wire FE_PHN2878_plain_text_43_;
   wire FE_PHN2877_plain_text_134_;
   wire FE_PHN2876_plain_text_13_;
   wire FE_PHN2875_plain_text_36_;
   wire FE_PHN2874_plain_text_26_;
   wire FE_PHN2873_n554;
   wire FE_PHN2872_n680;
   wire FE_PHN2871_plain_text_19_;
   wire FE_PHN2870_plain_text_239_;
   wire FE_PHN2869_n551;
   wire FE_PHN2868_plain_text_140_;
   wire FE_PHN2867_plain_text_50_;
   wire FE_PHN2866_n669;
   wire FE_PHN2865_plain_text_62_;
   wire FE_PHN2864_n756;
   wire FE_PHN2863_plain_text_130_;
   wire FE_PHN2862_plain_text_143_;
   wire FE_PHN2861_plain_text_64_;
   wire FE_PHN2860_plain_text_20_;
   wire FE_PHN2859_n651;
   wire FE_PHN2858_n636;
   wire FE_PHN2857_plain_text_197_;
   wire FE_PHN2854_n739;
   wire FE_PHN2853_n674;
   wire FE_PHN2852_n561;
   wire FE_PHN2851_n711;
   wire FE_PHN2822_plain_text_125_;
   wire FE_PHN2819_Din_127_;
   wire FE_PHN2818_Din_126_;
   wire FE_PHN2817_Din_31_;
   wire FE_PHN2815_n426;
   wire FE_PHN2804_pbv1;
   wire FE_PHN2801_pf0;
   wire FE_PHN2800_pbv0;
   wire FE_PHN2796_n385;
   wire FE_PHN2794_n474;
   wire FE_PHN2037_plain_text_124_;
   wire FE_PHN2035_plain_text_235_;
   wire FE_PHN2034_plain_text_154_;
   wire FE_PHN2033_plain_text_238_;
   wire FE_PHN2032_plain_text_226_;
   wire FE_PHN2031_plain_text_232_;
   wire FE_PHN2030_plain_text_219_;
   wire FE_PHN2029_plain_text_153_;
   wire FE_PHN2028_plain_text_172_;
   wire FE_PHN2027_plain_text_184_;
   wire FE_PHN2026_plain_text_209_;
   wire FE_PHN2025_plain_text_144_;
   wire FE_PHN2024_plain_text_165_;
   wire FE_PHN2023_plain_text_185_;
   wire FE_PHN2022_plain_text_38_;
   wire FE_PHN2021_plain_text_229_;
   wire FE_PHN2020_plain_text_242_;
   wire FE_PHN2019_plain_text_160_;
   wire FE_PHN2018_plain_text_204_;
   wire FE_PHN2017_plain_text_41_;
   wire FE_PHN2016_plain_text_35_;
   wire FE_PHN2015_plain_text_67_;
   wire FE_PHN2014_plain_text_195_;
   wire FE_PHN2013_plain_text_135_;
   wire FE_PHN2012_plain_text_233_;
   wire FE_PHN2011_plain_text_199_;
   wire FE_PHN2010_plain_text_245_;
   wire FE_PHN1999_Din_112_;
   wire FE_PHN1996_Din_4_;
   wire FE_PHN1995_Din_118_;
   wire FE_PHN1994_Din_113_;
   wire FE_PHN1993_Din_19_;
   wire FE_PHN1990_Din_119_;
   wire FE_PHN1988_Din_11_;
   wire FE_PHN1987_Din_17_;
   wire FE_PHN1986_Din_111_;
   wire FE_PHN1985_Din_115_;
   wire FE_PHN1984_Din_110_;
   wire FE_PHN1983_Din_13_;
   wire FE_PHN1982_Din_20_;
   wire FE_PHN1981_Din_105_;
   wire FE_PHN1980_Din_15_;
   wire FE_PHN1979_Din_18_;
   wire FE_PHN1978_Din_51_;
   wire FE_PHN1977_Din_54_;
   wire FE_PHN1976_Din_16_;
   wire FE_PHN1975_Din_85_;
   wire FE_PHN1973_Din_116_;
   wire FE_PHN1971_Din_100_;
   wire FE_PHN1970_Din_53_;
   wire FE_PHN1968_Din_83_;
   wire FE_PHN1967_Din_107_;
   wire FE_PHN1966_Din_87_;
   wire FE_PHN1964_Din_101_;
   wire FE_PHN1963_Din_86_;
   wire FE_PHN1961_Din_69_;
   wire FE_PHN1960_Din_52_;
   wire FE_PHN1956_Din_84_;
   wire FE_PHN1955_Din_108_;
   wire FE_PHN1954_Din_10_;
   wire FE_PHN1953_Din_77_;
   wire FE_PHN1952_Din_70_;
   wire FE_PHN1951_Din_102_;
   wire FE_PHN1950_Din_117_;
   wire FE_PHN1949_n615;
   wire FE_PHN1948_Din_109_;
   wire FE_PHN1947_n591;
   wire FE_PHN1946_n517;
   wire FE_PHN1945_Din_46_;
   wire FE_PHN1944_n691;
   wire FE_PHN1943_Din_78_;
   wire FE_PHN1942_Din_37_;
   wire FE_PHN1941_Din_45_;
   wire FE_PHN1940_Din_43_;
   wire FE_PHN1939_n687;
   wire FE_PHN1938_n528;
   wire FE_PHN1937_Din_97_;
   wire FE_PHN1936_n619;
   wire FE_PHN1935_n387;
   wire FE_PHN1934_n660;
   wire FE_PHN1933_n523;
   wire FE_PHN1932_n526;
   wire FE_PHN1931_n555;
   wire FE_PHN1929_n635;
   wire FE_PHN1928_n613;
   wire FE_PHN1927_n678;
   wire FE_PHN1926_n634;
   wire FE_PHN1925_Din_103_;
   wire FE_PHN1924_n560;
   wire FE_PHN1923_n618;
   wire FE_PHN1922_n559;
   wire FE_PHN1921_n755;
   wire FE_PHN1920_n583;
   wire FE_PHN1919_n556;
   wire FE_PHN1918_n649;
   wire FE_PHN1916_Din_99_;
   wire FE_PHN1915_n573;
   wire FE_PHN1914_n653;
   wire FE_PHN1913_Din_75_;
   wire FE_PHN1912_n527;
   wire FE_PHN1911_n735;
   wire FE_PHN1910_Din_104_;
   wire FE_PHN1909_n592;
   wire FE_PHN1908_Din_82_;
   wire FE_PHN1907_Din_76_;
   wire FE_PHN1906_n315;
   wire FE_PHN1904_n283;
   wire FE_PHN1903_n518;
   wire FE_PHN1902_n552;
   wire FE_PHN1901_n281;
   wire FE_PHN1900_n529;
   wire FE_PHN1898_n734;
   wire FE_PHN1897_n291;
   wire FE_PHN1896_Din_96_;
   wire FE_PHN1895_n692;
   wire FE_PHN1890_n549;
   wire FE_PHN1886_n524;
   wire FE_PHN1875_n581;
   wire FE_PHN1865_n679;
   wire FE_PHN1845_n553;
   wire FE_PHN1842_n616;
   wire FE_PHN1838_plain_text_248_;
   wire FE_PHN1836_n550;
   wire FE_PHN1825_n498;
   wire FE_PHN1815_n580;
   wire FE_PHN1753_n574;
   wire FE_PHN1741_n677;
   wire FE_PHN1704_n676;
   wire FE_PHN1465_n747;
   wire FE_PHN1462_plain_text_1_;
   wire FE_PHN1461_plain_text_0_;
   wire FE_PHN1460_plain_text_2_;
   wire FE_PHN1459_Din_120_;
   wire FE_PHN1453_plain_text_5_;
   wire FE_PHN1452_plain_text_123_;
   wire FE_PHN1451_plain_text_14_;
   wire FE_PHN1450_plain_text_6_;
   wire FE_PHN1448_plain_text_7_;
   wire FE_PHN1447_plain_text_214_;
   wire FE_PHN1443_plain_text_182_;
   wire FE_PHN1440_plain_text_132_;
   wire FE_PHN1439_plain_text_183_;
   wire FE_PHN1438_plain_text_122_;
   wire FE_PHN1437_n443;
   wire FE_PHN1436_plain_text_126_;
   wire FE_PHN1435_n386;
   wire FE_PHN1433_plain_text_246_;
   wire FE_PHN1432_plain_text_215_;
   wire FE_PHN1431_n475;
   wire FE_PHN1430_plain_text_179_;
   wire FE_PHN1428_plain_text_69_;
   wire FE_PHN1427_plain_text_147_;
   wire FE_PHN1426_plain_text_25_;
   wire FE_PHN1424_plain_text_12_;
   wire FE_PHN1423_n272;
   wire FE_PHN1420_plain_text_189_;
   wire FE_PHN1418_plain_text_205_;
   wire FE_PHN1417_plain_text_187_;
   wire FE_PHN1411_plain_text_171_;
   wire FE_PHN1410_plain_text_28_;
   wire FE_PHN1409_plain_text_210_;
   wire FE_PHN1407_n486;
   wire FE_PHN1403_plain_text_174_;
   wire FE_PHN1400_plain_text_240_;
   wire FE_PHN1399_plain_text_138_;
   wire FE_PHN1398_plain_text_228_;
   wire FE_PHN1396_plain_text_145_;
   wire FE_PHN1390_plain_text_178_;
   wire FE_PHN1389_plain_text_218_;
   wire FE_PHN1387_plain_text_139_;
   wire FE_PHN1386_plain_text_200_;
   wire FE_PHN1385_plain_text_177_;
   wire FE_PHN1384_plain_text_58_;
   wire FE_PHN1383_plain_text_18_;
   wire FE_PHN1382_plain_text_48_;
   wire FE_PHN1381_plain_text_216_;
   wire FE_PHN1379_plain_text_163_;
   wire FE_PHN1378_plain_text_196_;
   wire FE_PHN1377_plain_text_30_;
   wire FE_PHN1376_plain_text_194_;
   wire FE_PHN1374_plain_text_231_;
   wire FE_PHN1373_plain_text_202_;
   wire FE_PHN1372_plain_text_206_;
   wire FE_PHN1371_plain_text_169_;
   wire FE_PHN1370_plain_text_40_;
   wire FE_PHN1369_plain_text_65_;
   wire FE_PHN1368_plain_text_224_;
   wire FE_PHN1366_plain_text_114_;
   wire FE_PHN1365_plain_text_170_;
   wire FE_PHN1364_plain_text_136_;
   wire FE_PHN1363_plain_text_175_;
   wire FE_PHN1362_plain_text_72_;
   wire FE_PHN1361_plain_text_243_;
   wire FE_PHN1359_plain_text_42_;
   wire FE_PHN1358_plain_text_198_;
   wire FE_PHN1357_n423;
   wire FE_PHN1356_n456;
   wire FE_PHN1355_plain_text_32_;
   wire FE_PHN1354_plain_text_98_;
   wire FE_PHN1352_plain_text_79_;
   wire FE_PHN1351_plain_text_213_;
   wire FE_PHN1350_plain_text_176_;
   wire FE_PHN1349_plain_text_71_;
   wire FE_PHN1348_plain_text_80_;
   wire FE_PHN1347_plain_text_129_;
   wire FE_PHN1346_plain_text_230_;
   wire FE_PHN1344_plain_text_73_;
   wire FE_PHN1343_plain_text_81_;
   wire FE_PHN1342_plain_text_74_;
   wire FE_PHN1341_plain_text_142_;
   wire FE_PHN1340_n721;
   wire FE_PHN1339_plain_text_236_;
   wire FE_PHN1338_plain_text_50_;
   wire FE_PHN1337_plain_text_128_;
   wire FE_PHN1336_plain_text_239_;
   wire FE_PHN1334_plain_text_47_;
   wire FE_PHN1332_plain_text_44_;
   wire FE_PHN1331_plain_text_244_;
   wire FE_PHN1330_n425;
   wire FE_PHN1329_plain_text_201_;
   wire FE_PHN1328_plain_text_106_;
   wire FE_PHN1327_plain_text_141_;
   wire FE_PHN1325_plain_text_137_;
   wire FE_PHN1320_plain_text_68_;
   wire FE_PHN1319_n508;
   wire FE_PHN1317_plain_text_64_;
   wire FE_PHN1316_plain_text_34_;
   wire FE_PHN1309_Din_5_;
   wire FE_PHN1308_Din_2_;
   wire FE_PHN1307_Din_1_;
   wire FE_PHN1306_Din_38_;
   wire FE_PHN1305_Din_3_;
   wire FE_PHN1304_Din_0_;
   wire FE_PHN1303_Din_36_;
   wire FE_PHN1302_Din_7_;
   wire FE_PHN1301_Din_67_;
   wire FE_PHN1300_Din_68_;
   wire FE_PHN1298_Din_35_;
   wire FE_PHN1297_Din_71_;
   wire FE_PHN1296_Din_66_;
   wire FE_PHN1295_Din_6_;
   wire FE_PHN1294_Din_44_;
   wire FE_PHN1293_Din_64_;
   wire FE_PHN1292_Din_48_;
   wire FE_PHN1291_Din_80_;
   wire FE_PHN1290_Din_73_;
   wire FE_PHN1287_Din_74_;
   wire FE_PHN1286_Din_50_;
   wire FE_PHN1285_Din_40_;
   wire FE_PHN1283_Din_65_;
   wire FE_PHN1282_Din_106_;
   wire FE_PHN1281_Din_81_;
   wire FE_PHN1280_Din_42_;
   wire FE_PHN1279_Din_22_;
   wire FE_PHN1278_Din_114_;
   wire FE_PHN1277_Din_39_;
   wire FE_PHN1276_Din_79_;
   wire FE_PHN1275_Din_49_;
   wire FE_PHN1274_Din_98_;
   wire FE_PHN1273_Din_41_;
   wire FE_PHN1272_Din_9_;
   wire FE_PHN1271_Din_34_;
   wire FE_PHN1270_Din_32_;
   wire FE_PHN1269_Din_14_;
   wire FE_PHN1268_Din_8_;
   wire FE_PHN1267_Din_47_;
   wire FE_PHN1266_Din_72_;
   wire FE_PHN1260_Din_33_;
   wire FE_PHN1250_plain_text_251_;
   wire FE_PHN1248_plain_text_254_;
   wire FE_PHN1243_n812;
   wire FE_PHN1242_plain_text_250_;
   wire FE_PHN1240_plain_text_252_;
   wire FE_PHN1228_plain_text_253_;
   wire FE_PHN1218_plain_text_249_;
   wire FE_PHN1217_Din_121_;
   wire FE_PHN1216_Din_27_;
   wire FE_PHN1215_Din_28_;
   wire FE_PHN1214_Din_29_;
   wire FE_PHN1213_Din_123_;
   wire FE_PHN1212_n659;
   wire FE_PHN1210_plain_text_3_;
   wire FE_PHN1209_plain_text_157_;
   wire FE_PHN1208_plain_text_133_;
   wire FE_PHN1207_plain_text_118_;
   wire FE_PHN1206_plain_text_116_;
   wire FE_PHN1205_plain_text_24_;
   wire FE_PHN1204_plain_text_59_;
   wire FE_PHN1203_n546;
   wire FE_PHN1202_plain_text_17_;
   wire FE_PHN1201_plain_text_8_;
   wire FE_PHN1200_plain_text_109_;
   wire FE_PHN1199_plain_text_127_;
   wire FE_PHN1198_n625;
   wire FE_PHN1196_plain_text_54_;
   wire FE_PHN1195_plain_text_162_;
   wire FE_PHN1194_plain_text_152_;
   wire FE_PHN1193_plain_text_101_;
   wire FE_PHN1192_plain_text_22_;
   wire FE_PHN1191_plain_text_150_;
   wire FE_PHN1190_plain_text_146_;
   wire FE_PHN1189_plain_text_70_;
   wire FE_PHN1188_plain_text_121_;
   wire FE_PHN1187_plain_text_61_;
   wire FE_PHN1186_n609;
   wire FE_PHN1185_plain_text_186_;
   wire FE_PHN1184_plain_text_92_;
   wire FE_PHN1183_plain_text_223_;
   wire FE_PHN1182_plain_text_91_;
   wire FE_PHN1181_plain_text_78_;
   wire FE_PHN1180_plain_text_203_;
   wire FE_PHN1179_plain_text_208_;
   wire FE_PHN1178_plain_text_85_;
   wire FE_PHN1177_plain_text_112_;
   wire FE_PHN1176_plain_text_60_;
   wire FE_PHN1175_plain_text_99_;
   wire FE_PHN1174_plain_text_159_;
   wire FE_PHN1173_plain_text_117_;
   wire FE_PHN1171_plain_text_86_;
   wire FE_PHN1170_plain_text_11_;
   wire FE_PHN1169_plain_text_181_;
   wire FE_PHN1168_plain_text_173_;
   wire FE_PHN1167_plain_text_93_;
   wire FE_PHN1166_plain_text_16_;
   wire FE_PHN1165_plain_text_190_;
   wire FE_PHN1163_plain_text_168_;
   wire FE_PHN1162_plain_text_149_;
   wire FE_PHN1161_plain_text_193_;
   wire FE_PHN1160_plain_text_156_;
   wire FE_PHN1159_plain_text_37_;
   wire FE_PHN1158_plain_text_36_;
   wire FE_PHN1157_plain_text_29_;
   wire FE_PHN1156_plain_text_134_;
   wire FE_PHN1155_plain_text_9_;
   wire FE_PHN1154_n459;
   wire FE_PHN1153_plain_text_95_;
   wire FE_PHN1152_plain_text_158_;
   wire FE_PHN1151_plain_text_107_;
   wire FE_PHN1150_plain_text_19_;
   wire FE_PHN1149_plain_text_45_;
   wire FE_PHN1148_plain_text_120_;
   wire FE_PHN1147_plain_text_241_;
   wire FE_PHN1146_plain_text_83_;
   wire FE_PHN1145_plain_text_115_;
   wire FE_PHN1144_plain_text_131_;
   wire FE_PHN1143_plain_text_88_;
   wire FE_PHN1142_plain_text_89_;
   wire FE_PHN1141_plain_text_90_;
   wire FE_PHN1140_n710;
   wire FE_PHN1139_plain_text_234_;
   wire FE_PHN1138_plain_text_55_;
   wire FE_PHN1137_plain_text_222_;
   wire FE_PHN1136_n395;
   wire FE_PHN1135_plain_text_102_;
   wire FE_PHN1134_plain_text_148_;
   wire FE_PHN1133_plain_text_21_;
   wire FE_PHN1132_plain_text_207_;
   wire FE_PHN1131_plain_text_63_;
   wire FE_PHN1130_plain_text_221_;
   wire FE_PHN1129_plain_text_62_;
   wire FE_PHN1128_n434;
   wire FE_PHN1127_plain_text_161_;
   wire FE_PHN1126_plain_text_31_;
   wire FE_PHN1125_plain_text_23_;
   wire FE_PHN1124_plain_text_130_;
   wire FE_PHN1123_plain_text_110_;
   wire FE_PHN1122_plain_text_56_;
   wire FE_PHN1121_n725;
   wire FE_PHN1120_plain_text_108_;
   wire FE_PHN1119_plain_text_84_;
   wire FE_PHN1118_plain_text_211_;
   wire FE_PHN1117_plain_text_225_;
   wire FE_PHN1116_plain_text_97_;
   wire FE_PHN1115_plain_text_113_;
   wire FE_PHN1114_plain_text_66_;
   wire FE_PHN1113_plain_text_100_;
   wire FE_PHN1112_plain_text_104_;
   wire FE_PHN1111_plain_text_57_;
   wire FE_PHN1110_plain_text_103_;
   wire FE_PHN1109_plain_text_96_;
   wire FE_PHN1108_plain_text_192_;
   wire FE_PHN1106_plain_text_151_;
   wire FE_PHN1105_plain_text_220_;
   wire FE_PHN1104_plain_text_119_;
   wire FE_PHN1103_plain_text_76_;
   wire FE_PHN1102_plain_text_164_;
   wire FE_PHN1101_plain_text_87_;
   wire FE_PHN1099_plain_text_217_;
   wire FE_PHN1097_plain_text_82_;
   wire FE_PHN1095_plain_text_94_;
   wire FE_PHN1094_plain_text_143_;
   wire FE_PHN1091_plain_text_27_;
   wire FE_PHN1090_n639;
   wire FE_PHN1089_plain_text_49_;
   wire FE_PHN1082_plain_text_33_;
   wire FE_PHN1078_plain_text_105_;
   wire FE_PHN1073_plain_text_52_;
   wire FE_PHN1072_n668;
   wire FE_PHN1071_plain_text_111_;
   wire FE_PHN1070_n740;
   wire FE_PHN1069_plain_text_247_;
   wire FE_PHN1068_plain_text_51_;
   wire FE_PHN1065_plain_text_167_;
   wire FE_PHN1061_n644;
   wire FE_PHN1059_plain_text_188_;
   wire FE_PHN1047_plain_text_39_;
   wire FE_PHN1042_plain_text_53_;
   wire FE_PHN1039_plain_text_166_;
   wire FE_PHN911_Din_93_;
   wire FE_PHN910_Din_24_;
   wire FE_PHN909_Din_124_;
   wire FE_PHN908_Din_26_;
   wire FE_PHN907_Din_25_;
   wire FE_PHN906_Din_94_;
   wire FE_PHN904_Din_88_;
   wire FE_PHN903_Din_56_;
   wire FE_PHN902_Din_122_;
   wire FE_PHN901_Din_59_;
   wire FE_PHN900_Din_91_;
   wire FE_PHN899_Din_60_;
   wire FE_PHN898_Din_57_;
   wire FE_PHN897_Din_90_;
   wire FE_PHN895_Din_63_;
   wire FE_PHN894_Din_62_;
   wire FE_PHN893_Din_58_;
   wire FE_PHN892_Din_61_;
   wire FE_PHN891_Din_95_;
   wire FE_PHN890_Din_89_;
   wire FE_PHN889_Din_92_;
   wire FE_PHN888_plain_text_4_;
   wire FE_PHN886_plain_text_227_;
   wire FE_PHN884_plain_text_15_;
   wire FE_PHN883_plain_text_77_;
   wire FE_PHN882_plain_text_155_;
   wire FE_PHN880_plain_text_10_;
   wire FE_PHN875_plain_text_26_;
   wire FE_PHN874_plain_text_13_;
   wire FE_PHN870_plain_text_140_;
   wire FE_PHN864_plain_text_43_;
   wire FE_PHN861_plain_text_75_;
   wire FE_PHN860_plain_text_212_;
   wire FE_PHN837_plain_text_20_;
   wire FE_PHN835_plain_text_237_;
   wire FE_PHN830_plain_text_180_;
   wire FE_PHN829_plain_text_197_;
   wire FE_PHN828_plain_text_46_;
   wire FE_PHN824_plain_text_191_;
   wire FE_PHN823_n718;
   wire FE_PHN749_Din_125_;
   wire FE_PHN742_Din_30_;
   wire FE_PHN711_n427;
   wire FE_PHN704_n258;
   wire FE_PHN680_Din_183_;
   wire FE_PHN679_Din_182_;
   wire FE_PHN677_Din_158_;
   wire FE_PHN676_Din_157_;
   wire FE_PHN675_Din_155_;
   wire FE_PHN674_Din_147_;
   wire FE_PHN673_Din_148_;
   wire FE_PHN672_Din_156_;
   wire FE_PHN671_Din_149_;
   wire FE_PHN670_Din_211_;
   wire FE_PHN669_Din_146_;
   wire FE_PHN668_Din_186_;
   wire FE_PHN667_Din_159_;
   wire FE_PHN666_Din_180_;
   wire FE_PHN665_Din_188_;
   wire FE_PHN664_Din_250_;
   wire FE_PHN663_Din_225_;
   wire FE_PHN662_Din_208_;
   wire FE_PHN661_Din_181_;
   wire FE_PHN660_Din_151_;
   wire FE_PHN659_Din_247_;
   wire FE_PHN658_Din_252_;
   wire FE_PHN657_Din_212_;
   wire FE_PHN656_Din_150_;
   wire FE_PHN655_Din_140_;
   wire FE_PHN654_Din_220_;
   wire FE_PHN653_Din_227_;
   wire FE_PHN652_Din_237_;
   wire FE_PHN651_Din_221_;
   wire FE_PHN650_Din_249_;
   wire FE_PHN649_Din_244_;
   wire FE_PHN648_Din_241_;
   wire FE_PHN647_Din_255_;
   wire FE_PHN645_Din_251_;
   wire FE_PHN644_Din_166_;
   wire FE_PHN643_Din_164_;
   wire FE_PHN642_Din_253_;
   wire FE_PHN641_Din_191_;
   wire FE_PHN640_Din_254_;
   wire FE_PHN639_Din_197_;
   wire FE_PHN637_Din_167_;
   wire FE_PHN532_Din_219_;
   wire FE_PHN531_Din_139_;
   wire FE_PHN530_Din_154_;
   wire FE_PHN529_Din_189_;
   wire FE_PHN527_Din_187_;
   wire FE_PHN526_Din_210_;
   wire FE_PHN525_Din_202_;
   wire FE_PHN524_Din_228_;
   wire FE_PHN523_Din_160_;
   wire FE_PHN522_Din_246_;
   wire FE_PHN521_Din_130_;
   wire FE_PHN520_Din_226_;
   wire FE_PHN519_Din_185_;
   wire FE_PHN518_Din_153_;
   wire FE_PHN517_Din_236_;
   wire FE_PHN516_Din_231_;
   wire FE_PHN515_Din_134_;
   wire FE_PHN514_Din_218_;
   wire FE_PHN513_Din_203_;
   wire FE_PHN512_Din_200_;
   wire FE_PHN511_Din_141_;
   wire FE_PHN510_Din_177_;
   wire FE_PHN509_Din_204_;
   wire FE_PHN508_Din_195_;
   wire FE_PHN507_Din_213_;
   wire FE_PHN506_Din_178_;
   wire FE_PHN504_Din_179_;
   wire FE_PHN503_Din_142_;
   wire FE_PHN502_Din_184_;
   wire FE_PHN501_Din_222_;
   wire FE_PHN500_Din_217_;
   wire FE_PHN499_Din_229_;
   wire FE_PHN498_Din_233_;
   wire FE_PHN497_Din_205_;
   wire FE_PHN496_Din_173_;
   wire FE_PHN495_Din_162_;
   wire FE_PHN494_Din_196_;
   wire FE_PHN493_Din_163_;
   wire FE_PHN492_Din_224_;
   wire FE_PHN491_Din_152_;
   wire FE_PHN490_Din_234_;
   wire FE_PHN489_Din_199_;
   wire FE_PHN488_Din_168_;
   wire FE_PHN487_Din_194_;
   wire FE_PHN486_Din_243_;
   wire FE_PHN485_Din_176_;
   wire FE_PHN484_Din_169_;
   wire FE_PHN483_Din_230_;
   wire FE_PHN482_Din_135_;
   wire FE_PHN481_Din_190_;
   wire FE_PHN480_Din_239_;
   wire FE_PHN479_Din_193_;
   wire FE_PHN478_Din_192_;
   wire FE_PHN477_Din_235_;
   wire FE_PHN476_Din_245_;
   wire FE_PHN475_Din_223_;
   wire FE_PHN474_Din_242_;
   wire FE_PHN473_Din_138_;
   wire FE_PHN472_Din_174_;
   wire FE_PHN471_Din_145_;
   wire FE_PHN470_Din_206_;
   wire FE_PHN469_Din_207_;
   wire FE_PHN468_Din_171_;
   wire FE_PHN467_Din_201_;
   wire FE_PHN466_Din_144_;
   wire FE_PHN465_Din_165_;
   wire FE_PHN464_Din_216_;
   wire FE_PHN463_Din_170_;
   wire FE_PHN462_Din_128_;
   wire FE_PHN461_Din_136_;
   wire FE_PHN460_Din_143_;
   wire FE_PHN459_Din_238_;
   wire FE_PHN458_Din_131_;
   wire FE_PHN457_Din_129_;
   wire FE_PHN456_Din_232_;
   wire FE_PHN455_Din_209_;
   wire FE_PHN454_Din_198_;
   wire FE_PHN453_Din_240_;
   wire FE_PHN452_Din_172_;
   wire FE_PHN451_Din_133_;
   wire FE_PHN450_Din_161_;
   wire FE_PHN449_Din_132_;
   wire FE_PHN448_Din_137_;
   wire FE_PHN447_Din_175_;
   wire FE_PHN446_Din_248_;
   wire FE_PHN119_n1;
   wire FE_OFN75_n1;
   wire FE_OFN74_n1;
   wire FE_OFN73_n1;
   wire FE_OFN72_n1;
   wire FE_OFN71_n1;
   wire FE_OFN70_n1;
   wire FE_OFN69_n1;
   wire FE_OFN68_n1;
   wire FE_OFN67_n1;
   wire FE_OFN66_n258;
   wire FE_OFN65_n258;
   wire FE_OFN64_n258;
   wire FE_OFN63_n210;
   wire FE_OFN62_n210;
   wire FE_OFN61_n210;
   wire FE_OFN60_n210;
   wire FE_OFN59_n210;
   wire FE_OFN52_reset_n;
   wire pbv1;
   wire pbv0;
   wire pf1;
   wire pf0;
   wire n1;
   wire n258;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire n478;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire n556;
   wire n557;
   wire n558;
   wire n559;
   wire n560;
   wire n561;
   wire n562;
   wire n563;
   wire n564;
   wire n565;
   wire n566;
   wire n567;
   wire n568;
   wire n569;
   wire n570;
   wire n571;
   wire n572;
   wire n573;
   wire n574;
   wire n575;
   wire n576;
   wire n577;
   wire n578;
   wire n579;
   wire n580;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire n593;
   wire n594;
   wire n595;
   wire n596;
   wire n597;
   wire n598;
   wire n599;
   wire n600;
   wire n601;
   wire n602;
   wire n603;
   wire n604;
   wire n605;
   wire n606;
   wire n607;
   wire n608;
   wire n609;
   wire n610;
   wire n611;
   wire n612;
   wire n613;
   wire n614;
   wire n615;
   wire n616;
   wire n617;
   wire n618;
   wire n619;
   wire n620;
   wire n621;
   wire n622;
   wire n623;
   wire n624;
   wire n625;
   wire n626;
   wire n627;
   wire n628;
   wire n629;
   wire n630;
   wire n631;
   wire n632;
   wire n633;
   wire n634;
   wire n635;
   wire n636;
   wire n637;
   wire n638;
   wire n639;
   wire n640;
   wire n641;
   wire n642;
   wire n643;
   wire n644;
   wire n645;
   wire n646;
   wire n647;
   wire n648;
   wire n649;
   wire n650;
   wire n651;
   wire n652;
   wire n653;
   wire n654;
   wire n655;
   wire n656;
   wire n657;
   wire n658;
   wire n659;
   wire n660;
   wire n661;
   wire n662;
   wire n663;
   wire n664;
   wire n665;
   wire n666;
   wire n667;
   wire n668;
   wire n669;
   wire n670;
   wire n671;
   wire n672;
   wire n673;
   wire n674;
   wire n675;
   wire n676;
   wire n677;
   wire n678;
   wire n679;
   wire n680;
   wire n681;
   wire n682;
   wire n683;
   wire n684;
   wire n685;
   wire n686;
   wire n687;
   wire n688;
   wire n689;
   wire n690;
   wire n691;
   wire n692;
   wire n693;
   wire n694;
   wire n695;
   wire n696;
   wire n697;
   wire n698;
   wire n699;
   wire n700;
   wire n701;
   wire n702;
   wire n703;
   wire n704;
   wire n705;
   wire n706;
   wire n707;
   wire n708;
   wire n709;
   wire n710;
   wire n711;
   wire n712;
   wire n713;
   wire n714;
   wire n715;
   wire n716;
   wire n717;
   wire n718;
   wire n719;
   wire n720;
   wire n721;
   wire n722;
   wire n723;
   wire n724;
   wire n725;
   wire n726;
   wire n727;
   wire n728;
   wire n729;
   wire n730;
   wire n731;
   wire n732;
   wire n733;
   wire n734;
   wire n735;
   wire n736;
   wire n737;
   wire n738;
   wire n739;
   wire n740;
   wire n741;
   wire n742;
   wire n743;
   wire n744;
   wire n745;
   wire n746;
   wire n747;
   wire n748;
   wire n749;
   wire n750;
   wire n751;
   wire n752;
   wire n753;
   wire n754;
   wire n755;
   wire n756;
   wire n757;
   wire n758;
   wire n759;
   wire n760;
   wire n761;
   wire n762;
   wire n763;
   wire n764;
   wire n765;
   wire n766;
   wire n767;
   wire n768;
   wire n769;
   wire n770;
   wire n771;
   wire n52;
   wire n78;
   wire n153;
   wire n171;
   wire n210;
   wire n781;
   wire n782;
   wire n783;
   wire n784;
   wire n785;
   wire n786;
   wire n787;
   wire n788;
   wire n789;
   wire n790;
   wire n791;
   wire n792;
   wire n793;
   wire n794;
   wire n795;
   wire n796;
   wire n797;
   wire n798;
   wire n799;
   wire n800;
   wire n801;
   wire n802;
   wire n803;
   wire n804;
   wire n805;
   wire n806;
   wire n807;
   wire n808;
   wire n809;
   wire n810;
   wire n811;
   wire n812;
   wire n813;
   wire n814;
   wire n815;
   wire n816;
   wire n817;
   wire n818;
   wire n819;
   wire n820;
   wire n821;
   wire n822;
   wire n823;
   wire n824;
   wire n825;
   wire n826;
   wire n827;
   wire n828;
   wire n829;
   wire n830;
   wire n831;
   wire n832;
   wire n833;
   wire n834;
   wire n835;
   wire n836;
   wire n837;
   wire n838;
   wire n839;
   wire n840;
   wire n841;
   wire n842;
   wire n843;
   wire n844;
   wire n845;
   wire n846;
   wire n847;
   wire n848;
   wire n849;
   wire n850;
   wire n851;
   wire n852;
   wire n853;
   wire n854;
   wire n855;
   wire n856;
   wire n857;
   wire n858;
   wire n859;
   wire n860;
   wire n861;
   wire n862;
   wire n863;
   wire n864;
   wire n865;
   wire n866;
   wire n867;
   wire n868;
   wire n869;
   wire n870;
   wire n871;
   wire n872;
   wire n873;
   wire n874;
   wire n875;
   wire n876;
   wire n877;
   wire n878;
   wire n879;
   wire n880;
   wire n881;
   wire n882;
   wire n883;
   wire n884;
   wire n885;
   wire n886;
   wire n887;
   wire n888;
   wire n889;
   wire n890;
   wire n891;
   wire n892;
   wire n893;
   wire n894;
   wire n895;
   wire n896;
   wire n897;
   wire n898;
   wire n899;
   wire n900;
   wire n901;
   wire n902;
   wire n903;
   wire n904;
   wire n905;
   wire n906;
   wire n907;
   wire n908;
   wire n909;
   wire n910;
   wire n911;
   wire n912;
   wire n913;
   wire n914;
   wire n915;
   wire n916;
   wire n917;
   wire n918;
   wire n919;
   wire n920;
   wire n921;
   wire n922;
   wire n923;
   wire n924;
   wire n925;
   wire n926;
   wire n927;
   wire n928;
   wire n929;
   wire n930;
   wire n931;
   wire n932;
   wire n933;
   wire n934;
   wire n935;
   wire n936;
   wire n937;
   wire n938;
   wire n939;
   wire n940;
   wire n941;
   wire n942;
   wire n943;
   wire n944;
   wire n945;
   wire n946;
   wire n947;
   wire n948;
   wire n949;
   wire n950;
   wire n951;
   wire n952;
   wire n953;
   wire n954;
   wire n955;
   wire n956;
   wire n957;
   wire n958;
   wire n959;
   wire n960;
   wire n961;
   wire n962;
   wire n963;
   wire n964;
   wire n965;
   wire n966;
   wire n967;
   wire n968;
   wire n969;
   wire n970;
   wire n971;
   wire n972;
   wire n973;
   wire n974;
   wire n975;
   wire n976;
   wire n977;
   wire n978;
   wire n979;
   wire n980;
   wire n981;
   wire n982;
   wire n983;
   wire n984;
   wire n985;
   wire n986;
   wire n987;
   wire n988;
   wire n989;
   wire n990;
   wire n991;
   wire n992;
   wire n993;
   wire n994;
   wire n995;
   wire n996;
   wire n997;
   wire n998;
   wire n999;
   wire n1000;
   wire n1001;
   wire n1002;
   wire n1003;
   wire n1004;
   wire n1005;
   wire n1006;
   wire n1007;
   wire n1008;
   wire n1009;
   wire n1010;
   wire n1011;
   wire n1012;
   wire n1013;
   wire n1014;
   wire n1015;
   wire n1016;
   wire n1017;
   wire n1018;
   wire n1019;
   wire n1020;
   wire n1021;
   wire n1022;
   wire n1023;
   wire n1024;
   wire n1025;
   wire n1026;
   wire n1027;
   wire n1028;
   wire n1029;
   wire n1030;
   wire n1031;
   wire n1032;
   wire n1033;
   wire n1034;
   wire n1035;
   wire n1036;
   wire [255:0] plain_text;

   BUFXL FE_PHC5257_plain_text_28_ (.Y(FE_PHN5257_plain_text_28_), 
	.A(FE_PHN3147_plain_text_28_));
   BUFXL FE_PHC5255_plain_text_185_ (.Y(FE_PHN5255_plain_text_185_), 
	.A(FE_PHN5240_plain_text_185_));
   CLKBUFX1 FE_PHC5254_n505 (.Y(FE_PHN5254_n505), 
	.A(FE_PHN5241_n505));
   BUFXL FE_PHC5243_plain_text_78_ (.Y(FE_PHN5243_plain_text_78_), 
	.A(plain_text[78]));
   BUFXL FE_PHC5242_plain_text_12_ (.Y(FE_PHN5242_plain_text_12_), 
	.A(FE_PHN3559_plain_text_12_));
   CLKBUFX1 FE_PHC5241_n505 (.Y(FE_PHN5241_n505), 
	.A(n505));
   CLKBUFX3 FE_PHC5240_plain_text_185_ (.Y(FE_PHN5240_plain_text_185_), 
	.A(plain_text[185]));
   DLY1X1 FE_PHC5239_plain_text_153_ (.Y(FE_PHN5239_plain_text_153_), 
	.A(plain_text[153]));
   DLY2X1 FE_PHC5238_n484 (.Y(FE_PHN5238_n484), 
	.A(n484));
   DLY2X1 FE_PHC5237_n420 (.Y(FE_PHN5237_n420), 
	.A(n420));
   DLY3X1 FE_PHC5236_plain_text_106_ (.Y(FE_PHN5236_plain_text_106_), 
	.A(plain_text[106]));
   BUFXL FE_PHC5234_plain_text_121_ (.Y(FE_PHN5234_plain_text_121_), 
	.A(FE_PHN3016_plain_text_121_));
   DLY2X1 FE_PHC5232_n516 (.Y(FE_PHN5232_n516), 
	.A(FE_PHN5157_n516));
   DLY2X1 FE_PHC5231_plain_text_49_ (.Y(FE_PHN5231_plain_text_49_), 
	.A(FE_PHN5156_plain_text_49_));
   BUFXL FE_PHC5230_Din_241_ (.Y(FE_PHN5230_Din_241_), 
	.A(FE_PHN648_Din_241_));
   BUFXL FE_PHC5171_plain_text_49_ (.Y(FE_PHN5171_plain_text_49_), 
	.A(FE_PHN5231_plain_text_49_));
   BUFXL FE_PHC5170_plain_text_1_ (.Y(FE_PHN5170_plain_text_1_), 
	.A(FE_PHN5155_plain_text_1_));
   BUFXL FE_PHC5158_n502 (.Y(FE_PHN5158_n502), 
	.A(FE_PHN3024_n502));
   CLKBUFX1 FE_PHC5157_n516 (.Y(FE_PHN5157_n516), 
	.A(FE_PHN2879_n516));
   CLKBUFX3 FE_PHC5156_plain_text_49_ (.Y(FE_PHN5156_plain_text_49_), 
	.A(plain_text[49]));
   CLKBUFX3 FE_PHC5155_plain_text_1_ (.Y(FE_PHN5155_plain_text_1_), 
	.A(FE_PHN3182_plain_text_1_));
   DLY2X1 FE_PHC5154_plain_text_121_ (.Y(FE_PHN5154_plain_text_121_), 
	.A(plain_text[121]));
   BUFXL FE_PHC5072_plain_text_125_ (.Y(FE_PHN5072_plain_text_125_), 
	.A(FE_PHN2822_plain_text_125_));
   DLY4X1 FE_PHC5069_pf0 (.Y(FE_PHN5069_pf0), 
	.A(FE_PHN2801_pf0));
   DLY4X1 FE_PHC5067_pbv0 (.Y(FE_PHN5067_pbv0), 
	.A(FE_PHN2800_pbv0));
   DLY2X1 FE_PHC5048_n475 (.Y(FE_PHN5048_n475), 
	.A(n475));
   DLY2X1 FE_PHC5046_n474 (.Y(FE_PHN5046_n474), 
	.A(n474));
   DLY2X1 FE_PHC3610_n265 (.Y(FE_PHN3610_n265), 
	.A(n265));
   DLY2X1 FE_PHC3609_n383 (.Y(FE_PHN3609_n383), 
	.A(n383));
   DLY2X1 FE_PHC3608_n262 (.Y(FE_PHN3608_n262), 
	.A(n262));
   DLY4X1 FE_PHC3607_plain_text_235_ (.Y(FE_PHN3607_plain_text_235_), 
	.A(plain_text[235]));
   DLY4X1 FE_PHC3606_n261 (.Y(FE_PHN3606_n261), 
	.A(n261));
   DLY3X1 FE_PHC3605_n285 (.Y(FE_PHN3605_n285), 
	.A(n285));
   DLY3X1 FE_PHC3604_n399 (.Y(FE_PHN3604_n399), 
	.A(n399));
   DLY4X1 FE_PHC3603_n442 (.Y(FE_PHN3603_n442), 
	.A(n442));
   DLY3X1 FE_PHC3602_n417 (.Y(FE_PHN3602_n417), 
	.A(n417));
   DLY3X1 FE_PHC3601_n382 (.Y(FE_PHN3601_n382), 
	.A(n382));
   DLY4X1 FE_PHC3600_n407 (.Y(FE_PHN3600_n407), 
	.A(n407));
   DLY3X1 FE_PHC3599_n329 (.Y(FE_PHN3599_n329), 
	.A(n329));
   DLY4X1 FE_PHC3598_n470 (.Y(FE_PHN3598_n470), 
	.A(n470));
   DLY4X1 FE_PHC3597_plain_text_172_ (.Y(FE_PHN3597_plain_text_172_), 
	.A(plain_text[172]));
   DLY3X1 FE_PHC3596_n270 (.Y(FE_PHN3596_n270), 
	.A(n270));
   DLY3X1 FE_PHC3595_n278 (.Y(FE_PHN3595_n278), 
	.A(n278));
   DLY4X1 FE_PHC3594_n284 (.Y(FE_PHN3594_n284), 
	.A(n284));
   DLY4X1 FE_PHC3593_n271 (.Y(FE_PHN3593_n271), 
	.A(n271));
   DLY3X1 FE_PHC3592_n267 (.Y(FE_PHN3592_n267), 
	.A(n267));
   DLY4X1 FE_PHC3591_n277 (.Y(FE_PHN3591_n277), 
	.A(n277));
   DLY4X1 FE_PHC3590_n409 (.Y(FE_PHN3590_n409), 
	.A(n409));
   DLY3X1 FE_PHC3589_n260 (.Y(FE_PHN3589_n260), 
	.A(n260));
   DLY4X1 FE_PHC3588_plain_text_204_ (.Y(FE_PHN3588_plain_text_204_), 
	.A(FE_PHN2018_plain_text_204_));
   DLY3X1 FE_PHC3587_n319 (.Y(FE_PHN3587_n319), 
	.A(n319));
   DLY4X1 FE_PHC3586_n264 (.Y(FE_PHN3586_n264), 
	.A(n264));
   DLY3X1 FE_PHC3585_n318 (.Y(FE_PHN3585_n318), 
	.A(n318));
   DLY3X1 FE_PHC3584_n263 (.Y(FE_PHN3584_n263), 
	.A(n263));
   DLY3X1 FE_PHC3583_n314 (.Y(FE_PHN3583_n314), 
	.A(n314));
   DLY4X1 FE_PHC3582_n488 (.Y(FE_PHN3582_n488), 
	.A(n488));
   DLY3X1 FE_PHC3581_n351 (.Y(FE_PHN3581_n351), 
	.A(n351));
   DLY3X1 FE_PHC3580_n506 (.Y(FE_PHN3580_n506), 
	.A(n506));
   DLY4X1 FE_PHC3579_n367 (.Y(FE_PHN3579_n367), 
	.A(n367));
   DLY4X1 FE_PHC3578_n266 (.Y(FE_PHN3578_n266), 
	.A(n266));
   DLY4X1 FE_PHC3577_n288 (.Y(FE_PHN3577_n288), 
	.A(n288));
   DLY3X1 FE_PHC3576_plain_text_139_ (.Y(FE_PHN3576_plain_text_139_), 
	.A(FE_PHN1387_plain_text_139_));
   DLY3X1 FE_PHC3575_n378 (.Y(FE_PHN3575_n378), 
	.A(n378));
   DLY3X1 FE_PHC3574_n472 (.Y(FE_PHN3574_n472), 
	.A(n472));
   DLY3X1 FE_PHC3573_n372 (.Y(FE_PHN3573_n372), 
	.A(n372));
   DLY4X1 FE_PHC3572_n374 (.Y(FE_PHN3572_n374), 
	.A(n374));
   DLY4X1 FE_PHC3571_n448 (.Y(FE_PHN3571_n448), 
	.A(n448));
   DLY4X1 FE_PHC3570_n415 (.Y(FE_PHN3570_n415), 
	.A(n415));
   DLY4X1 FE_PHC3569_n381 (.Y(FE_PHN3569_n381), 
	.A(n381));
   DLY4X1 FE_PHC3568_n449 (.Y(FE_PHN3568_n449), 
	.A(n449));
   DLY3X1 FE_PHC3567_n295 (.Y(FE_PHN3567_n295), 
	.A(n295));
   DLY3X1 FE_PHC3566_n331 (.Y(FE_PHN3566_n331), 
	.A(n331));
   DLY3X1 FE_PHC3565_n316 (.Y(FE_PHN3565_n316), 
	.A(n316));
   DLY3X1 FE_PHC3564_n333 (.Y(FE_PHN3564_n333), 
	.A(n333));
   DLY4X1 FE_PHC3563_n353 (.Y(FE_PHN3563_n353), 
	.A(n353));
   DLY4X1 FE_PHC3562_n274 (.Y(FE_PHN3562_n274), 
	.A(n274));
   DLY4X1 FE_PHC3561_n462 (.Y(FE_PHN3561_n462), 
	.A(n462));
   DLY4X1 FE_PHC3560_n380 (.Y(FE_PHN3560_n380), 
	.A(n380));
   DLY3X1 FE_PHC3559_plain_text_12_ (.Y(FE_PHN3559_plain_text_12_), 
	.A(FE_PHN1424_plain_text_12_));
   DLY3X1 FE_PHC3558_n439 (.Y(FE_PHN3558_n439), 
	.A(n439));
   DLY4X1 FE_PHC3557_n328 (.Y(FE_PHN3557_n328), 
	.A(n328));
   DLY4X1 FE_PHC3556_n317 (.Y(FE_PHN3556_n317), 
	.A(n317));
   DLY4X1 FE_PHC3555_n406 (.Y(FE_PHN3555_n406), 
	.A(n406));
   DLY4X1 FE_PHC3554_n468 (.Y(FE_PHN3554_n468), 
	.A(n468));
   DLY3X1 FE_PHC3553_n369 (.Y(FE_PHN3553_n369), 
	.A(n369));
   DLY3X1 FE_PHC3552_n273 (.Y(FE_PHN3552_n273), 
	.A(n273));
   DLY3X1 FE_PHC3551_n289 (.Y(FE_PHN3551_n289), 
	.A(n289));
   DLY3X1 FE_PHC3550_n401 (.Y(FE_PHN3550_n401), 
	.A(n401));
   DLY3X1 FE_PHC3549_n416 (.Y(FE_PHN3549_n416), 
	.A(n416));
   DLY4X1 FE_PHC3548_n339 (.Y(FE_PHN3548_n339), 
	.A(n339));
   DLY4X1 FE_PHC3547_n363 (.Y(FE_PHN3547_n363), 
	.A(n363));
   DLY3X1 FE_PHC3546_n345 (.Y(FE_PHN3546_n345), 
	.A(n345));
   DLY3X1 FE_PHC3545_n460 (.Y(FE_PHN3545_n460), 
	.A(n460));
   DLY3X1 FE_PHC3544_n446 (.Y(FE_PHN3544_n446), 
	.A(n446));
   DLY3X1 FE_PHC3543_n300 (.Y(FE_PHN3543_n300), 
	.A(n300));
   DLY3X1 FE_PHC3542_n355 (.Y(FE_PHN3542_n355), 
	.A(n355));
   DLY4X1 FE_PHC3541_n365 (.Y(FE_PHN3541_n365), 
	.A(n365));
   DLY4X1 FE_PHC3540_n361 (.Y(FE_PHN3540_n361), 
	.A(n361));
   DLY4X1 FE_PHC3539_n438 (.Y(FE_PHN3539_n438), 
	.A(n438));
   DLY4X1 FE_PHC3538_n349 (.Y(FE_PHN3538_n349), 
	.A(n349));
   DLY4X1 FE_PHC3537_n390 (.Y(FE_PHN3537_n390), 
	.A(n390));
   DLY4X1 FE_PHC3536_n292 (.Y(FE_PHN3536_n292), 
	.A(n292));
   DLY3X1 FE_PHC3535_n275 (.Y(FE_PHN3535_n275), 
	.A(n275));
   DLY3X1 FE_PHC3534_n463 (.Y(FE_PHN3534_n463), 
	.A(n463));
   DLY3X1 FE_PHC3533_n330 (.Y(FE_PHN3533_n330), 
	.A(n330));
   DLY3X1 FE_PHC3532_n337 (.Y(FE_PHN3532_n337), 
	.A(n337));
   DLY3X1 FE_PHC3531_n375 (.Y(FE_PHN3531_n375), 
	.A(n375));
   DLY4X1 FE_PHC3530_n282 (.Y(FE_PHN3530_n282), 
	.A(n282));
   DLY4X1 FE_PHC3529_n394 (.Y(FE_PHN3529_n394), 
	.A(n394));
   DLY4X1 FE_PHC3528_n308 (.Y(FE_PHN3528_n308), 
	.A(n308));
   DLY4X1 FE_PHC3527_n326 (.Y(FE_PHN3527_n326), 
	.A(n326));
   DLY4X1 FE_PHC3526_n366 (.Y(FE_PHN3526_n366), 
	.A(n366));
   DLY4X1 FE_PHC3525_n344 (.Y(FE_PHN3525_n344), 
	.A(n344));
   DLY4X1 FE_PHC3524_n352 (.Y(FE_PHN3524_n352), 
	.A(n352));
   DLY4X1 FE_PHC3523_n362 (.Y(FE_PHN3523_n362), 
	.A(n362));
   DLY4X1 FE_PHC3522_n307 (.Y(FE_PHN3522_n307), 
	.A(n307));
   DLY3X1 FE_PHC3521_n342 (.Y(FE_PHN3521_n342), 
	.A(n342));
   DLY3X1 FE_PHC3520_n303 (.Y(FE_PHN3520_n303), 
	.A(n303));
   DLY3X1 FE_PHC3519_n348 (.Y(FE_PHN3519_n348), 
	.A(n348));
   DLY3X1 FE_PHC3518_n485 (.Y(FE_PHN3518_n485), 
	.A(n485));
   DLY3X1 FE_PHC3517_n503 (.Y(FE_PHN3517_n503), 
	.A(n503));
   DLY4X1 FE_PHC3516_n371 (.Y(FE_PHN3516_n371), 
	.A(n371));
   DLY4X1 FE_PHC3515_n296 (.Y(FE_PHN3515_n296), 
	.A(n296));
   DLY4X1 FE_PHC3514_n477 (.Y(FE_PHN3514_n477), 
	.A(n477));
   DLY4X1 FE_PHC3513_n405 (.Y(FE_PHN3513_n405), 
	.A(n405));
   DLY3X1 FE_PHC3512_n334 (.Y(FE_PHN3512_n334), 
	.A(n334));
   DLY3X1 FE_PHC3511_n433 (.Y(FE_PHN3511_n433), 
	.A(n433));
   DLY3X1 FE_PHC3510_n357 (.Y(FE_PHN3510_n357), 
	.A(n357));
   DLY3X1 FE_PHC3509_n321 (.Y(FE_PHN3509_n321), 
	.A(n321));
   DLY3X1 FE_PHC3508_n441 (.Y(FE_PHN3508_n441), 
	.A(n441));
   DLY3X1 FE_PHC3507_n276 (.Y(FE_PHN3507_n276), 
	.A(n276));
   DLY3X1 FE_PHC3506_n400 (.Y(FE_PHN3506_n400), 
	.A(n400));
   DLY3X1 FE_PHC3505_n341 (.Y(FE_PHN3505_n341), 
	.A(n341));
   DLY3X1 FE_PHC3504_n496 (.Y(FE_PHN3504_n496), 
	.A(n496));
   DLY4X1 FE_PHC3503_n354 (.Y(FE_PHN3503_n354), 
	.A(n354));
   DLY4X1 FE_PHC3502_n280 (.Y(FE_PHN3502_n280), 
	.A(n280));
   DLY4X1 FE_PHC3501_n324 (.Y(FE_PHN3501_n324), 
	.A(n324));
   DLY4X1 FE_PHC3500_n379 (.Y(FE_PHN3500_n379), 
	.A(n379));
   DLY4X1 FE_PHC3499_n454 (.Y(FE_PHN3499_n454), 
	.A(n454));
   DLY3X1 FE_PHC3498_n482 (.Y(FE_PHN3498_n482), 
	.A(n482));
   DLY3X1 FE_PHC3497_n480 (.Y(FE_PHN3497_n480), 
	.A(n480));
   DLY3X1 FE_PHC3496_n325 (.Y(FE_PHN3496_n325), 
	.A(n325));
   DLY3X1 FE_PHC3495_n450 (.Y(FE_PHN3495_n450), 
	.A(n450));
   DLY4X1 FE_PHC3494_n473 (.Y(FE_PHN3494_n473), 
	.A(n473));
   DLY4X1 FE_PHC3493_n452 (.Y(FE_PHN3493_n452), 
	.A(n452));
   DLY4X1 FE_PHC3492_n440 (.Y(FE_PHN3492_n440), 
	.A(n440));
   DLY4X1 FE_PHC3491_n320 (.Y(FE_PHN3491_n320), 
	.A(n320));
   DLY4X1 FE_PHC3490_n279 (.Y(FE_PHN3490_n279), 
	.A(n279));
   DLY4X1 FE_PHC3489_n286 (.Y(FE_PHN3489_n286), 
	.A(n286));
   DLY3X1 FE_PHC3488_n297 (.Y(FE_PHN3488_n297), 
	.A(n297));
   DLY3X1 FE_PHC3487_n364 (.Y(FE_PHN3487_n364), 
	.A(n364));
   DLY3X1 FE_PHC3486_n350 (.Y(FE_PHN3486_n350), 
	.A(n350));
   DLY4X1 FE_PHC3485_n310 (.Y(FE_PHN3485_n310), 
	.A(n310));
   DLY4X1 FE_PHC3484_n347 (.Y(FE_PHN3484_n347), 
	.A(n347));
   DLY4X1 FE_PHC3483_n359 (.Y(FE_PHN3483_n359), 
	.A(n359));
   DLY4X1 FE_PHC3482_n312 (.Y(FE_PHN3482_n312), 
	.A(n312));
   DLY4X1 FE_PHC3481_n304 (.Y(FE_PHN3481_n304), 
	.A(n304));
   DLY4X1 FE_PHC3480_n302 (.Y(FE_PHN3480_n302), 
	.A(n302));
   DLY3X1 FE_PHC3479_n343 (.Y(FE_PHN3479_n343), 
	.A(n343));
   DLY3X1 FE_PHC3478_n465 (.Y(FE_PHN3478_n465), 
	.A(n465));
   DLY3X1 FE_PHC3477_n311 (.Y(FE_PHN3477_n311), 
	.A(n311));
   DLY3X1 FE_PHC3476_n346 (.Y(FE_PHN3476_n346), 
	.A(n346));
   DLY3X1 FE_PHC3475_n293 (.Y(FE_PHN3475_n293), 
	.A(n293));
   DLY4X1 FE_PHC3474_n306 (.Y(FE_PHN3474_n306), 
	.A(n306));
   DLY3X1 FE_PHC3473_n338 (.Y(FE_PHN3473_n338), 
	.A(n338));
   DLY4X1 FE_PHC3472_n373 (.Y(FE_PHN3472_n373), 
	.A(n373));
   DLY4X1 FE_PHC3471_n428 (.Y(FE_PHN3471_n428), 
	.A(n428));
   DLY4X1 FE_PHC3470_n499 (.Y(FE_PHN3470_n499), 
	.A(n499));
   DLY4X1 FE_PHC3469_n269 (.Y(FE_PHN3469_n269), 
	.A(n269));
   DLY3X1 FE_PHC3468_n429 (.Y(FE_PHN3468_n429), 
	.A(n429));
   DLY3X1 FE_PHC3467_n309 (.Y(FE_PHN3467_n309), 
	.A(n309));
   DLY4X1 FE_PHC3466_n393 (.Y(FE_PHN3466_n393), 
	.A(n393));
   DLY3X1 FE_PHC3465_n340 (.Y(FE_PHN3465_n340), 
	.A(n340));
   DLY4X1 FE_PHC3464_n268 (.Y(FE_PHN3464_n268), 
	.A(n268));
   DLY4X1 FE_PHC3463_n305 (.Y(FE_PHN3463_n305), 
	.A(n305));
   DLY4X1 FE_PHC3462_n476 (.Y(FE_PHN3462_n476), 
	.A(n476));
   DLY4X1 FE_PHC3461_n335 (.Y(FE_PHN3461_n335), 
	.A(n335));
   DLY4X1 FE_PHC3460_n421 (.Y(FE_PHN3460_n421), 
	.A(n421));
   DLY4X1 FE_PHC3459_n368 (.Y(FE_PHN3459_n368), 
	.A(n368));
   DLY4X1 FE_PHC3458_n356 (.Y(FE_PHN3458_n356), 
	.A(n356));
   DLY4X1 FE_PHC3457_n389 (.Y(FE_PHN3457_n389), 
	.A(n389));
   DLY3X1 FE_PHC3456_n332 (.Y(FE_PHN3456_n332), 
	.A(n332));
   DLY4X1 FE_PHC3455_n453 (.Y(FE_PHN3455_n453), 
	.A(n453));
   DLY4X1 FE_PHC3454_n392 (.Y(FE_PHN3454_n392), 
	.A(n392));
   DLY4X1 FE_PHC3453_n322 (.Y(FE_PHN3453_n322), 
	.A(n322));
   DLY4X1 FE_PHC3452_n294 (.Y(FE_PHN3452_n294), 
	.A(n294));
   DLY3X1 FE_PHC3451_n391 (.Y(FE_PHN3451_n391), 
	.A(n391));
   DLY4X1 FE_PHC3450_n336 (.Y(FE_PHN3450_n336), 
	.A(n336));
   DLY4X1 FE_PHC3449_n358 (.Y(FE_PHN3449_n358), 
	.A(n358));
   DLY4X1 FE_PHC3448_n388 (.Y(FE_PHN3448_n388), 
	.A(n388));
   DLY4X1 FE_PHC3447_n403 (.Y(FE_PHN3447_n403), 
	.A(n403));
   DLY3X1 FE_PHC3446_n360 (.Y(FE_PHN3446_n360), 
	.A(n360));
   DLY4X1 FE_PHC3445_n500 (.Y(FE_PHN3445_n500), 
	.A(n500));
   DLY4X1 FE_PHC3443_n483 (.Y(FE_PHN3443_n483), 
	.A(n483));
   DLY4X1 FE_PHC3442_n398 (.Y(FE_PHN3442_n398), 
	.A(n398));
   DLY4X1 FE_PHC3441_n431 (.Y(FE_PHN3441_n431), 
	.A(n431));
   DLY4X1 FE_PHC3440_n430 (.Y(FE_PHN3440_n430), 
	.A(n430));
   DLY3X1 FE_PHC3439_n461 (.Y(FE_PHN3439_n461), 
	.A(n461));
   DLY4X1 FE_PHC3438_n299 (.Y(FE_PHN3438_n299), 
	.A(n299));
   DLY4X1 FE_PHC3436_n397 (.Y(FE_PHN3436_n397), 
	.A(n397));
   DLY3X1 FE_PHC3432_n313 (.Y(FE_PHN3432_n313), 
	.A(n313));
   DLY4X1 FE_PHC3405_n491 (.Y(FE_PHN3405_n491), 
	.A(n491));
   DLY4X1 FE_PHC3404_plain_text_32_ (.Y(FE_PHN3404_plain_text_32_), 
	.A(plain_text[32]));
   DLY3X1 FE_PHC3402_n410 (.Y(FE_PHN3402_n410), 
	.A(n410));
   DLY3X1 FE_PHC3401_n419 (.Y(FE_PHN3401_n419), 
	.A(n419));
   DLY4X1 FE_PHC3400_plain_text_42_ (.Y(FE_PHN3400_plain_text_42_), 
	.A(plain_text[42]));
   DLY3X1 FE_PHC3399_n418 (.Y(FE_PHN3399_n418), 
	.A(n418));
   DLY4X1 FE_PHC3398_n323 (.Y(FE_PHN3398_n323), 
	.A(n323));
   DLY4X1 FE_PHC3397_n467 (.Y(FE_PHN3397_n467), 
	.A(n467));
   DLY4X1 FE_PHC3396_n411 (.Y(FE_PHN3396_n411), 
	.A(n411));
   DLY4X1 FE_PHC3395_n466 (.Y(FE_PHN3395_n466), 
	.A(n466));
   DLY3X1 FE_PHC3394_n490 (.Y(FE_PHN3394_n490), 
	.A(n490));
   DLY4X1 FE_PHC3393_n435 (.Y(FE_PHN3393_n435), 
	.A(n435));
   DLY3X1 FE_PHC3392_n458 (.Y(FE_PHN3392_n458), 
	.A(n458));
   DLY2X1 FE_PHC3391_plain_text_0_ (.Y(FE_PHN3391_plain_text_0_), 
	.A(FE_PHN1461_plain_text_0_));
   DLY4X1 FE_PHC3390_plain_text_147_ (.Y(FE_PHN3390_plain_text_147_), 
	.A(plain_text[147]));
   DLY4X1 FE_PHC3389_plain_text_157_ (.Y(FE_PHN3389_plain_text_157_), 
	.A(FE_PHN1209_plain_text_157_));
   DLY4X1 FE_PHC3387_n624 (.Y(FE_PHN3387_n624), 
	.A(n624));
   DLY4X1 FE_PHC3386_plain_text_133_ (.Y(FE_PHN3386_plain_text_133_), 
	.A(FE_PHN1208_plain_text_133_));
   DLY4X1 FE_PHC3385_n620 (.Y(FE_PHN3385_n620), 
	.A(n620));
   DLY4X1 FE_PHC3384_n709 (.Y(FE_PHN3384_n709), 
	.A(n709));
   DLY4X1 FE_PHC3383_n724 (.Y(FE_PHN3383_n724), 
	.A(n724));
   DLY3X1 FE_PHC3382_plain_text_18_ (.Y(FE_PHN3382_plain_text_18_), 
	.A(FE_PHN1383_plain_text_18_));
   DLY3X1 FE_PHC3381_n686 (.Y(FE_PHN3381_n686), 
	.A(n686));
   DLY4X1 FE_PHC3380_n638 (.Y(FE_PHN3380_n638), 
	.A(n638));
   DLY3X1 FE_PHC3379_plain_text_33_ (.Y(FE_PHN3379_plain_text_33_), 
	.A(plain_text[33]));
   DLY3X1 FE_PHC3377_n542 (.Y(FE_PHN3377_n542), 
	.A(n542));
   DLY3X1 FE_PHC3376_plain_text_59_ (.Y(FE_PHN3376_plain_text_59_), 
	.A(FE_PHN1204_plain_text_59_));
   DLY3X1 FE_PHC3375_n545 (.Y(FE_PHN3375_n545), 
	.A(n545));
   DLY3X1 FE_PHC3374_n584 (.Y(FE_PHN3374_n584), 
	.A(n584));
   DLY3X1 FE_PHC3372_n543 (.Y(FE_PHN3372_n543), 
	.A(n543));
   DLY3X1 FE_PHC3370_n658 (.Y(FE_PHN3370_n658), 
	.A(n658));
   DLY3X1 FE_PHC3369_plain_text_146_ (.Y(FE_PHN3369_plain_text_146_), 
	.A(FE_PHN1190_plain_text_146_));
   DLY3X1 FE_PHC3368_n608 (.Y(FE_PHN3368_n608), 
	.A(n608));
   DLY3X1 FE_PHC3367_plain_text_196_ (.Y(FE_PHN3367_plain_text_196_), 
	.A(FE_PHN1378_plain_text_196_));
   DLY3X1 FE_PHC3366_n605 (.Y(FE_PHN3366_n605), 
	.A(n605));
   DLY4X1 FE_PHC3364_n582 (.Y(FE_PHN3364_n582), 
	.A(n582));
   DLY4X1 FE_PHC3363_plain_text_163_ (.Y(FE_PHN3363_plain_text_163_), 
	.A(FE_PHN1379_plain_text_163_));
   DLY3X1 FE_PHC3361_n693 (.Y(FE_PHN3361_n693), 
	.A(n693));
   DLY4X1 FE_PHC3357_n519 (.Y(FE_PHN3357_n519), 
	.A(n519));
   DLY4X1 FE_PHC3355_plain_text_225_ (.Y(FE_PHN3355_plain_text_225_), 
	.A(FE_PHN1117_plain_text_225_));
   DLY4X1 FE_PHC3354_plain_text_168_ (.Y(FE_PHN3354_plain_text_168_), 
	.A(plain_text[168]));
   DLY3X1 FE_PHC3352_n617 (.Y(FE_PHN3352_n617), 
	.A(n617));
   DLY3X1 FE_PHC3350_plain_text_203_ (.Y(FE_PHN3350_plain_text_203_), 
	.A(plain_text[203]));
   DLY4X1 FE_PHC3348_plain_text_52_ (.Y(FE_PHN3348_plain_text_52_), 
	.A(plain_text[52]));
   DLY4X1 FE_PHC3347_n736 (.Y(FE_PHN3347_n736), 
	.A(n736));
   DLY3X1 FE_PHC3346_n557 (.Y(FE_PHN3346_n557), 
	.A(n557));
   DLY3X1 FE_PHC3337_plain_text_241_ (.Y(FE_PHN3337_plain_text_241_), 
	.A(plain_text[241]));
   DLY4X1 FE_PHC3336_plain_text_243_ (.Y(FE_PHN3336_plain_text_243_), 
	.A(FE_PHN1361_plain_text_243_));
   DLY3X1 FE_PHC3320_plain_text_55_ (.Y(FE_PHN3320_plain_text_55_), 
	.A(plain_text[55]));
   DLY3X1 FE_PHC3318_plain_text_23_ (.Y(FE_PHN3318_plain_text_23_), 
	.A(plain_text[23]));
   DLY4X1 FE_PHC3317_n768 (.Y(FE_PHN3317_n768), 
	.A(n768));
   DLY4X1 FE_PHC3311_plain_text_193_ (.Y(FE_PHN3311_plain_text_193_), 
	.A(FE_PHN1161_plain_text_193_));
   DLY3X1 FE_PHC3306_n726 (.Y(FE_PHN3306_n726), 
	.A(n726));
   DLY4X1 FE_PHC3300_n612 (.Y(FE_PHN3300_n612), 
	.A(n612));
   DLY4X1 FE_PHC3299_plain_text_31_ (.Y(FE_PHN3299_plain_text_31_), 
	.A(plain_text[31]));
   DLY4X1 FE_PHC3298_plain_text_161_ (.Y(FE_PHN3298_plain_text_161_), 
	.A(plain_text[161]));
   DLY4X1 FE_PHC3297_n558 (.Y(FE_PHN3297_n558), 
	.A(n558));
   DLY4X1 FE_PHC3291_n741 (.Y(FE_PHN3291_n741), 
	.A(n741));
   DLY4X1 FE_PHC3287_plain_text_192_ (.Y(FE_PHN3287_plain_text_192_), 
	.A(plain_text[192]));
   DLY4X1 FE_PHC3286_n522 (.Y(FE_PHN3286_n522), 
	.A(n522));
   DLY4X1 FE_PHC3280_plain_text_21_ (.Y(FE_PHN3280_plain_text_21_), 
	.A(plain_text[21]));
   DLY4X1 FE_PHC3279_n704 (.Y(FE_PHN3279_n704), 
	.A(n704));
   DLY4X1 FE_PHC3264_n645 (.Y(FE_PHN3264_n645), 
	.A(n645));
   DLY4X1 FE_PHC3257_n661 (.Y(FE_PHN3257_n661), 
	.A(n661));
   DLY4X1 FE_PHC3254_n765 (.Y(FE_PHN3254_n765), 
	.A(n765));
   DLY4X1 FE_PHC3199_n606 (.Y(FE_PHN3199_n606), 
	.A(n606));
   DLY2X1 FE_PHC3182_plain_text_1_ (.Y(FE_PHN3182_plain_text_1_), 
	.A(plain_text[1]));
   DLY2X1 FE_PHC3181_plain_text_2_ (.Y(FE_PHN3181_plain_text_2_), 
	.A(plain_text[2]));
   DLY3X1 FE_PHC3176_plain_text_123_ (.Y(FE_PHN3176_plain_text_123_), 
	.A(plain_text[123]));
   DLY4X1 FE_PHC3175_plain_text_6_ (.Y(FE_PHN3175_plain_text_6_), 
	.A(plain_text[6]));
   DLY4X1 FE_PHC3174_plain_text_14_ (.Y(FE_PHN3174_plain_text_14_), 
	.A(FE_PHN1451_plain_text_14_));
   DLY4X1 FE_PHC3172_n717 (.Y(FE_PHN3172_n717), 
	.A(n717));
   DLY3X1 FE_PHC3171_plain_text_7_ (.Y(FE_PHN3171_plain_text_7_), 
	.A(FE_PHN1448_plain_text_7_));
   DLY3X1 FE_PHC3170_n771 (.Y(FE_PHN3170_n771), 
	.A(n771));
   DLY4X1 FE_PHC3169_plain_text_182_ (.Y(FE_PHN3169_plain_text_182_), 
	.A(FE_PHN1443_plain_text_182_));
   DLY3X1 FE_PHC3168_n716 (.Y(FE_PHN3168_n716), 
	.A(n716));
   DLY4X1 FE_PHC3167_plain_text_122_ (.Y(FE_PHN3167_plain_text_122_), 
	.A(plain_text[122]));
   DLY4X1 FE_PHC3166_plain_text_179_ (.Y(FE_PHN3166_plain_text_179_), 
	.A(plain_text[179]));
   DLY3X1 FE_PHC3165_plain_text_25_ (.Y(FE_PHN3165_plain_text_25_), 
	.A(FE_PHN1426_plain_text_25_));
   DLY3X1 FE_PHC3164_plain_text_69_ (.Y(FE_PHN3164_plain_text_69_), 
	.A(FE_PHN1428_plain_text_69_));
   DLY4X1 FE_PHC3163_plain_text_11_ (.Y(FE_PHN3163_plain_text_11_), 
	.A(plain_text[11]));
   DLY3X1 FE_PHC3162_plain_text_228_ (.Y(FE_PHN3162_plain_text_228_), 
	.A(plain_text[228]));
   DLY4X1 FE_PHC3159_n744 (.Y(FE_PHN3159_n744), 
	.A(n744));
   DLY3X1 FE_PHC3158_n712 (.Y(FE_PHN3158_n712), 
	.A(n712));
   DLY4X1 FE_PHC3157_plain_text_231_ (.Y(FE_PHN3157_plain_text_231_), 
	.A(plain_text[231]));
   DLY3X1 FE_PHC3156_plain_text_171_ (.Y(FE_PHN3156_plain_text_171_), 
	.A(plain_text[171]));
   DLY4X1 FE_PHC3155_n723 (.Y(FE_PHN3155_n723), 
	.A(n723));
   DLY4X1 FE_PHC3154_plain_text_189_ (.Y(FE_PHN3154_plain_text_189_), 
	.A(FE_PHN1420_plain_text_189_));
   DLY4X1 FE_PHC3153_plain_text_205_ (.Y(FE_PHN3153_plain_text_205_), 
	.A(FE_PHN1418_plain_text_205_));
   DLY3X1 FE_PHC3152_plain_text_210_ (.Y(FE_PHN3152_plain_text_210_), 
	.A(FE_PHN1409_plain_text_210_));
   DLY3X1 FE_PHC3151_plain_text_48_ (.Y(FE_PHN3151_plain_text_48_), 
	.A(plain_text[48]));
   DLY4X1 FE_PHC3150_n746 (.Y(FE_PHN3150_n746), 
	.A(n746));
   DLY3X1 FE_PHC3148_plain_text_178_ (.Y(FE_PHN3148_plain_text_178_), 
	.A(FE_PHN1390_plain_text_178_));
   DLY3X1 FE_PHC3147_plain_text_28_ (.Y(FE_PHN3147_plain_text_28_), 
	.A(FE_PHN1410_plain_text_28_));
   DLY3X1 FE_PHC3146_plain_text_65_ (.Y(FE_PHN3146_plain_text_65_), 
	.A(plain_text[65]));
   DLY4X1 FE_PHC3145_n748 (.Y(FE_PHN3145_n748), 
	.A(n748));
   DLY3X1 FE_PHC3144_n713 (.Y(FE_PHN3144_n713), 
	.A(n713));
   DLY3X1 FE_PHC3143_plain_text_206_ (.Y(FE_PHN3143_plain_text_206_), 
	.A(FE_PHN1372_plain_text_206_));
   DLY3X1 FE_PHC3142_n641 (.Y(FE_PHN3142_n641), 
	.A(n641));
   DLY4X1 FE_PHC3141_plain_text_54_ (.Y(FE_PHN3141_plain_text_54_), 
	.A(plain_text[54]));
   DLY3X1 FE_PHC3140_n714 (.Y(FE_PHN3140_n714), 
	.A(n714));
   DLY3X1 FE_PHC3139_plain_text_198_ (.Y(FE_PHN3139_plain_text_198_), 
	.A(plain_text[198]));
   DLY3X1 FE_PHC3138_n715 (.Y(FE_PHN3138_n715), 
	.A(n715));
   DLY3X1 FE_PHC3137_plain_text_138_ (.Y(FE_PHN3137_plain_text_138_), 
	.A(FE_PHN1399_plain_text_138_));
   DLY4X1 FE_PHC3136_plain_text_216_ (.Y(FE_PHN3136_plain_text_216_), 
	.A(FE_PHN1381_plain_text_216_));
   DLY4X1 FE_PHC3135_plain_text_56_ (.Y(FE_PHN3135_plain_text_56_), 
	.A(plain_text[56]));
   DLY4X1 FE_PHC3134_n525 (.Y(FE_PHN3134_n525), 
	.A(n525));
   DLY3X1 FE_PHC3133_plain_text_170_ (.Y(FE_PHN3133_plain_text_170_), 
	.A(plain_text[170]));
   DLY4X1 FE_PHC3132_n539 (.Y(FE_PHN3132_n539), 
	.A(n539));
   DLY3X1 FE_PHC3131_plain_text_169_ (.Y(FE_PHN3131_plain_text_169_), 
	.A(FE_PHN1371_plain_text_169_));
   DLY4X1 FE_PHC3130_n745 (.Y(FE_PHN3130_n745), 
	.A(n745));
   DLY3X1 FE_PHC3129_n750 (.Y(FE_PHN3129_n750), 
	.A(n750));
   DLY3X1 FE_PHC3128_plain_text_81_ (.Y(FE_PHN3128_plain_text_81_), 
	.A(plain_text[81]));
   DLY4X1 FE_PHC3127_n754 (.Y(FE_PHN3127_n754), 
	.A(n754));
   DLY4X1 FE_PHC3126_plain_text_141_ (.Y(FE_PHN3126_plain_text_141_), 
	.A(plain_text[141]));
   DLY4X1 FE_PHC3125_plain_text_68_ (.Y(FE_PHN3125_plain_text_68_), 
	.A(plain_text[68]));
   DLY4X1 FE_PHC3124_plain_text_72_ (.Y(FE_PHN3124_plain_text_72_), 
	.A(FE_PHN1362_plain_text_72_));
   DLY4X1 FE_PHC3123_n537 (.Y(FE_PHN3123_n537), 
	.A(n537));
   DLY4X1 FE_PHC3122_n530 (.Y(FE_PHN3122_n530), 
	.A(n530));
   DLY4X1 FE_PHC3121_plain_text_128_ (.Y(FE_PHN3121_plain_text_128_), 
	.A(FE_PHN1337_plain_text_128_));
   DLY3X1 FE_PHC3120_n751 (.Y(FE_PHN3120_n751), 
	.A(n751));
   DLY4X1 FE_PHC3119_n743 (.Y(FE_PHN3119_n743), 
	.A(n743));
   DLY4X1 FE_PHC3118_n722 (.Y(FE_PHN3118_n722), 
	.A(n722));
   DLY4X1 FE_PHC3117_n749 (.Y(FE_PHN3117_n749), 
	.A(n749));
   DLY3X1 FE_PHC3116_plain_text_175_ (.Y(FE_PHN3116_plain_text_175_), 
	.A(FE_PHN1363_plain_text_175_));
   DLY4X1 FE_PHC3115_n719 (.Y(FE_PHN3115_n719), 
	.A(n719));
   DLY4X1 FE_PHC3114_plain_text_137_ (.Y(FE_PHN3114_plain_text_137_), 
	.A(plain_text[137]));
   DLY4X1 FE_PHC3113_n562 (.Y(FE_PHN3113_n562), 
	.A(n562));
   DLY4X1 FE_PHC3112_plain_text_129_ (.Y(FE_PHN3112_plain_text_129_), 
	.A(FE_PHN1347_plain_text_129_));
   DLY4X1 FE_PHC3111_n640 (.Y(FE_PHN3111_n640), 
	.A(n640));
   DLY4X1 FE_PHC3110_plain_text_47_ (.Y(FE_PHN3110_plain_text_47_), 
	.A(plain_text[47]));
   DLY4X1 FE_PHC3109_n538 (.Y(FE_PHN3109_n538), 
	.A(n538));
   DLY3X1 FE_PHC3103_plain_text_10_ (.Y(FE_PHN3103_plain_text_10_), 
	.A(FE_PHN880_plain_text_10_));
   DLY4X1 FE_PHC3102_plain_text_118_ (.Y(FE_PHN3102_plain_text_118_), 
	.A(FE_PHN1207_plain_text_118_));
   DLY4X1 FE_PHC3101_plain_text_227_ (.Y(FE_PHN3101_plain_text_227_), 
	.A(FE_PHN886_plain_text_227_));
   DLY3X1 FE_PHC3100_plain_text_212_ (.Y(FE_PHN3100_plain_text_212_), 
	.A(plain_text[212]));
   DLY4X1 FE_PHC3099_plain_text_162_ (.Y(FE_PHN3099_plain_text_162_), 
	.A(FE_PHN1195_plain_text_162_));
   DLY3X1 FE_PHC3098_plain_text_60_ (.Y(FE_PHN3098_plain_text_60_), 
	.A(plain_text[60]));
   DLY3X1 FE_PHC3097_plain_text_150_ (.Y(FE_PHN3097_plain_text_150_), 
	.A(FE_PHN1191_plain_text_150_));
   DLY4X1 FE_PHC3096_plain_text_234_ (.Y(FE_PHN3096_plain_text_234_), 
	.A(FE_PHN1139_plain_text_234_));
   DLY4X1 FE_PHC3093_plain_text_217_ (.Y(FE_PHN3093_plain_text_217_), 
	.A(plain_text[217]));
   DLY4X1 FE_PHC3092_plain_text_75_ (.Y(FE_PHN3092_plain_text_75_), 
	.A(FE_PHN861_plain_text_75_));
   DLY4X1 FE_PHC3090_plain_text_49_ (.Y(FE_PHN3090_plain_text_49_), 
	.A(FE_PHN5171_plain_text_49_));
   DLY4X1 FE_PHC3088_plain_text_251_ (.Y(FE_PHN3088_plain_text_251_), 
	.A(plain_text[251]));
   DLY4X1 FE_PHC3087_plain_text_254_ (.Y(FE_PHN3087_plain_text_254_), 
	.A(FE_PHN1248_plain_text_254_));
   DLY4X1 FE_PHC3086_plain_text_180_ (.Y(FE_PHN3086_plain_text_180_), 
	.A(plain_text[180]));
   DLY4X1 FE_PHC3084_plain_text_191_ (.Y(FE_PHN3084_plain_text_191_), 
	.A(FE_PHN824_plain_text_191_));
   DLY4X1 FE_PHC3083_plain_text_46_ (.Y(FE_PHN3083_plain_text_46_), 
	.A(plain_text[46]));
   DLY4X1 FE_PHC3082_plain_text_249_ (.Y(FE_PHN3082_plain_text_249_), 
	.A(plain_text[249]));
   DLY2X1 FE_PHC3080_n384 (.Y(FE_PHN3080_n384), 
	.A(n384));
   DLY3X1 FE_PHC3079_plain_text_5_ (.Y(FE_PHN3079_plain_text_5_), 
	.A(FE_PHN1453_plain_text_5_));
   DLY2X1 FE_PHC3078_n479 (.Y(FE_PHN3078_n479), 
	.A(n479));
   DLY4X1 FE_PHC3077_n414 (.Y(FE_PHN3077_n414), 
	.A(n414));
   DLY3X1 FE_PHC3076_n447 (.Y(FE_PHN3076_n447), 
	.A(n447));
   DLY4X1 FE_PHC3075_n298 (.Y(FE_PHN3075_n298), 
	.A(n298));
   DLY4X1 FE_PHC3074_plain_text_3_ (.Y(FE_PHN3074_plain_text_3_), 
	.A(plain_text[3]));
   DLY3X1 FE_PHC3073_n420 (.Y(FE_PHN3073_n420), 
	.A(FE_PHN5237_n420));
   DLY4X1 FE_PHC3072_n437 (.Y(FE_PHN3072_n437), 
	.A(n437));
   DLY4X1 FE_PHC3071_n478 (.Y(FE_PHN3071_n478), 
	.A(n478));
   DLY3X1 FE_PHC3070_n481 (.Y(FE_PHN3070_n481), 
	.A(n481));
   DLY3X1 FE_PHC3069_n445 (.Y(FE_PHN3069_n445), 
	.A(n445));
   DLY4X1 FE_PHC3068_n413 (.Y(FE_PHN3068_n413), 
	.A(n413));
   DLY4X1 FE_PHC3067_n376 (.Y(FE_PHN3067_n376), 
	.A(n376));
   DLY3X1 FE_PHC3066_n301 (.Y(FE_PHN3066_n301), 
	.A(n301));
   DLY4X1 FE_PHC3065_plain_text_246_ (.Y(FE_PHN3065_plain_text_246_), 
	.A(FE_PHN1433_plain_text_246_));
   DLY4X1 FE_PHC3064_n377 (.Y(FE_PHN3064_n377), 
	.A(n377));
   DLY4X1 FE_PHC3063_plain_text_58_ (.Y(FE_PHN3063_plain_text_58_), 
	.A(plain_text[58]));
   DLY4X1 FE_PHC3062_n412 (.Y(FE_PHN3062_n412), 
	.A(n412));
   DLY3X1 FE_PHC3061_n327 (.Y(FE_PHN3061_n327), 
	.A(n327));
   DLY3X1 FE_PHC3060_n464 (.Y(FE_PHN3060_n464), 
	.A(n464));
   DLY3X1 FE_PHC3059_n455 (.Y(FE_PHN3059_n455), 
	.A(n455));
   DLY4X1 FE_PHC3058_n436 (.Y(FE_PHN3058_n436), 
	.A(n436));
   DLY4X1 FE_PHC3057_n290 (.Y(FE_PHN3057_n290), 
	.A(n290));
   DLY4X1 FE_PHC3056_n487 (.Y(FE_PHN3056_n487), 
	.A(n487));
   DLY3X1 FE_PHC3055_n504 (.Y(FE_PHN3055_n504), 
	.A(n504));
   DLY3X1 FE_PHC3054_plain_text_24_ (.Y(FE_PHN3054_plain_text_24_), 
	.A(FE_PHN1205_plain_text_24_));
   DLY4X1 FE_PHC3053_n444 (.Y(FE_PHN3053_n444), 
	.A(n444));
   DLY3X1 FE_PHC3052_plain_text_114_ (.Y(FE_PHN3052_plain_text_114_), 
	.A(FE_PHN1366_plain_text_114_));
   DLY3X1 FE_PHC3051_plain_text_93_ (.Y(FE_PHN3051_plain_text_93_), 
	.A(plain_text[93]));
   DLY3X1 FE_PHC3050_n515 (.Y(FE_PHN3050_n515), 
	.A(n515));
   DLY3X1 FE_PHC3049_n497 (.Y(FE_PHN3049_n497), 
	.A(n497));
   DLY3X1 FE_PHC3048_plain_text_73_ (.Y(FE_PHN3048_plain_text_73_), 
	.A(plain_text[73]));
   DLY3X1 FE_PHC3047_n493 (.Y(FE_PHN3047_n493), 
	.A(n493));
   DLY4X1 FE_PHC3046_n484 (.Y(FE_PHN3046_n484), 
	.A(FE_PHN5238_n484));
   DLY3X1 FE_PHC3045_plain_text_190_ (.Y(FE_PHN3045_plain_text_190_), 
	.A(FE_PHN1165_plain_text_190_));
   DLY3X1 FE_PHC3044_plain_text_17_ (.Y(FE_PHN3044_plain_text_17_), 
	.A(FE_PHN1202_plain_text_17_));
   DLY3X1 FE_PHC3043_plain_text_109_ (.Y(FE_PHN3043_plain_text_109_), 
	.A(FE_PHN1200_plain_text_109_));
   DLY4X1 FE_PHC3042_n287 (.Y(FE_PHN3042_n287), 
	.A(n287));
   DLY4X1 FE_PHC3041_plain_text_95_ (.Y(FE_PHN3041_plain_text_95_), 
	.A(plain_text[95]));
   DLY3X1 FE_PHC3040_plain_text_200_ (.Y(FE_PHN3040_plain_text_200_), 
	.A(FE_PHN1386_plain_text_200_));
   DLY3X1 FE_PHC3039_n370 (.Y(FE_PHN3039_n370), 
	.A(n370));
   DLY4X1 FE_PHC3038_plain_text_101_ (.Y(FE_PHN3038_plain_text_101_), 
	.A(FE_PHN1193_plain_text_101_));
   DLY4X1 FE_PHC3037_plain_text_107_ (.Y(FE_PHN3037_plain_text_107_), 
	.A(FE_PHN1151_plain_text_107_));
   DLY4X1 FE_PHC3036_n489 (.Y(FE_PHN3036_n489), 
	.A(n489));
   DLY3X1 FE_PHC3035_n471 (.Y(FE_PHN3035_n471), 
	.A(n471));
   DLY3X1 FE_PHC3034_plain_text_29_ (.Y(FE_PHN3034_plain_text_29_), 
	.A(FE_PHN1157_plain_text_29_));
   DLY3X1 FE_PHC3033_plain_text_103_ (.Y(FE_PHN3033_plain_text_103_), 
	.A(plain_text[103]));
   DLY4X1 FE_PHC3032_plain_text_120_ (.Y(FE_PHN3032_plain_text_120_), 
	.A(plain_text[120]));
   DLY4X1 FE_PHC3031_plain_text_202_ (.Y(FE_PHN3031_plain_text_202_), 
	.A(FE_PHN1373_plain_text_202_));
   DLY4X1 FE_PHC3030_plain_text_112_ (.Y(FE_PHN3030_plain_text_112_), 
	.A(FE_PHN1177_plain_text_112_));
   DLY4X1 FE_PHC3029_plain_text_22_ (.Y(FE_PHN3029_plain_text_22_), 
	.A(FE_PHN1192_plain_text_22_));
   DLY4X1 FE_PHC3028_n422 (.Y(FE_PHN3028_n422), 
	.A(n422));
   DLY3X1 FE_PHC3027_plain_text_79_ (.Y(FE_PHN3027_plain_text_79_), 
	.A(FE_PHN1352_plain_text_79_));
   DLY3X1 FE_PHC3026_n505 (.Y(FE_PHN3026_n505), 
	.A(FE_PHN5254_n505));
   DLY3X1 FE_PHC3025_plain_text_131_ (.Y(FE_PHN3025_plain_text_131_), 
	.A(FE_PHN1144_plain_text_131_));
   DLY3X1 FE_PHC3024_n502 (.Y(FE_PHN3024_n502), 
	.A(n502));
   DLY4X1 FE_PHC3023_plain_text_207_ (.Y(FE_PHN3023_plain_text_207_), 
	.A(plain_text[207]));
   DLY4X1 FE_PHC3022_n402 (.Y(FE_PHN3022_n402), 
	.A(n402));
   DLY4X1 FE_PHC3021_n396 (.Y(FE_PHN3021_n396), 
	.A(n396));
   DLY3X1 FE_PHC3020_plain_text_99_ (.Y(FE_PHN3020_plain_text_99_), 
	.A(FE_PHN1175_plain_text_99_));
   DLY3X1 FE_PHC3019_plain_text_115_ (.Y(FE_PHN3019_plain_text_115_), 
	.A(plain_text[115]));
   DLY4X1 FE_PHC3018_n501 (.Y(FE_PHN3018_n501), 
	.A(n501));
   DLY3X1 FE_PHC3017_plain_text_90_ (.Y(FE_PHN3017_plain_text_90_), 
	.A(FE_PHN1141_plain_text_90_));
   DLY3X1 FE_PHC3016_plain_text_121_ (.Y(FE_PHN3016_plain_text_121_), 
	.A(FE_PHN1188_plain_text_121_));
   DLY4X1 FE_PHC3015_plain_text_91_ (.Y(FE_PHN3015_plain_text_91_), 
	.A(FE_PHN1182_plain_text_91_));
   DLY4X1 FE_PHC3014_n494 (.Y(FE_PHN3014_n494), 
	.A(n494));
   DLY4X1 FE_PHC3013_plain_text_70_ (.Y(FE_PHN3013_plain_text_70_), 
	.A(FE_PHN1189_plain_text_70_));
   DLY4X1 FE_PHC3012_plain_text_194_ (.Y(FE_PHN3012_plain_text_194_), 
	.A(FE_PHN1376_plain_text_194_));
   DLY4X1 FE_PHC3011_plain_text_61_ (.Y(FE_PHN3011_plain_text_61_), 
	.A(plain_text[61]));
   DLY4X1 FE_PHC3010_plain_text_149_ (.Y(FE_PHN3010_plain_text_149_), 
	.A(FE_PHN1162_plain_text_149_));
   DLY4X1 FE_PHC3009_plain_text_89_ (.Y(FE_PHN3009_plain_text_89_), 
	.A(plain_text[89]));
   DLY4X1 FE_PHC3008_plain_text_208_ (.Y(FE_PHN3008_plain_text_208_), 
	.A(FE_PHN1179_plain_text_208_));
   DLY4X1 FE_PHC3007_plain_text_156_ (.Y(FE_PHN3007_plain_text_156_), 
	.A(plain_text[156]));
   DLY4X1 FE_PHC3006_plain_text_84_ (.Y(FE_PHN3006_plain_text_84_), 
	.A(plain_text[84]));
   DLY3X1 FE_PHC3005_plain_text_66_ (.Y(FE_PHN3005_plain_text_66_), 
	.A(plain_text[66]));
   DLY3X1 FE_PHC3004_plain_text_223_ (.Y(FE_PHN3004_plain_text_223_), 
	.A(FE_PHN1183_plain_text_223_));
   DLY3X1 FE_PHC3003_plain_text_159_ (.Y(FE_PHN3003_plain_text_159_), 
	.A(FE_PHN1174_plain_text_159_));
   DLY3X1 FE_PHC3002_plain_text_71_ (.Y(FE_PHN3002_plain_text_71_), 
	.A(plain_text[71]));
   DLY3X1 FE_PHC3001_plain_text_82_ (.Y(FE_PHN3001_plain_text_82_), 
	.A(plain_text[82]));
   DLY3X1 FE_PHC3000_plain_text_78_ (.Y(FE_PHN3000_plain_text_78_), 
	.A(FE_PHN1181_plain_text_78_));
   DLY3X1 FE_PHC2999_plain_text_57_ (.Y(FE_PHN2999_plain_text_57_), 
	.A(plain_text[57]));
   DLY3X1 FE_PHC2998_plain_text_92_ (.Y(FE_PHN2998_plain_text_92_), 
	.A(FE_PHN1184_plain_text_92_));
   DLY3X1 FE_PHC2997_n495 (.Y(FE_PHN2997_n495), 
	.A(n495));
   DLY4X1 FE_PHC2996_n492 (.Y(FE_PHN2996_n492), 
	.A(n492));
   DLY3X1 FE_PHC2995_plain_text_85_ (.Y(FE_PHN2995_plain_text_85_), 
	.A(FE_PHN1178_plain_text_85_));
   DLY3X1 FE_PHC2994_plain_text_186_ (.Y(FE_PHN2994_plain_text_186_), 
	.A(FE_PHN1185_plain_text_186_));
   DLY4X1 FE_PHC2992_plain_text_98_ (.Y(FE_PHN2992_plain_text_98_), 
	.A(FE_PHN1354_plain_text_98_));
   DLY4X1 FE_PHC2991_plain_text_106_ (.Y(FE_PHN2991_plain_text_106_), 
	.A(FE_PHN1328_plain_text_106_));
   DLY4X1 FE_PHC2989_plain_text_181_ (.Y(FE_PHN2989_plain_text_181_), 
	.A(plain_text[181]));
   DLY3X1 FE_PHC2988_plain_text_173_ (.Y(FE_PHN2988_plain_text_173_), 
	.A(plain_text[173]));
   DLY3X1 FE_PHC2987_plain_text_86_ (.Y(FE_PHN2987_plain_text_86_), 
	.A(FE_PHN1171_plain_text_86_));
   DLY4X1 FE_PHC2986_n507 (.Y(FE_PHN2986_n507), 
	.A(n507));
   DLY4X1 FE_PHC2985_plain_text_74_ (.Y(FE_PHN2985_plain_text_74_), 
	.A(plain_text[74]));
   DLY4X1 FE_PHC2984_plain_text_158_ (.Y(FE_PHN2984_plain_text_158_), 
	.A(plain_text[158]));
   DLY4X1 FE_PHC2981_plain_text_102_ (.Y(FE_PHN2981_plain_text_102_), 
	.A(FE_PHN1135_plain_text_102_));
   DLY3X1 FE_PHC2980_plain_text_94_ (.Y(FE_PHN2980_plain_text_94_), 
	.A(plain_text[94]));
   DLY3X1 FE_PHC2979_plain_text_104_ (.Y(FE_PHN2979_plain_text_104_), 
	.A(plain_text[104]));
   DLY3X1 FE_PHC2978_plain_text_37_ (.Y(FE_PHN2978_plain_text_37_), 
	.A(FE_PHN1159_plain_text_37_));
   DLY3X1 FE_PHC2977_plain_text_80_ (.Y(FE_PHN2977_plain_text_80_), 
	.A(FE_PHN1348_plain_text_80_));
   DLY3X1 FE_PHC2976_plain_text_164_ (.Y(FE_PHN2976_plain_text_164_), 
	.A(plain_text[164]));
   DLY3X1 FE_PHC2975_n424 (.Y(FE_PHN2975_n424), 
	.A(n424));
   DLY4X1 FE_PHC2974_n404 (.Y(FE_PHN2974_n404), 
	.A(n404));
   DLY4X1 FE_PHC2973_plain_text_96_ (.Y(FE_PHN2973_plain_text_96_), 
	.A(FE_PHN1109_plain_text_96_));
   DLY4X1 FE_PHC2972_plain_text_87_ (.Y(FE_PHN2972_plain_text_87_), 
	.A(plain_text[87]));
   DLY4X1 FE_PHC2971_plain_text_9_ (.Y(FE_PHN2971_plain_text_9_), 
	.A(FE_PHN1155_plain_text_9_));
   DLY4X1 FE_PHC2969_plain_text_213_ (.Y(FE_PHN2969_plain_text_213_), 
	.A(FE_PHN1351_plain_text_213_));
   DLY4X1 FE_PHC2968_plain_text_220_ (.Y(FE_PHN2968_plain_text_220_), 
	.A(plain_text[220]));
   DLY4X1 FE_PHC2967_n432 (.Y(FE_PHN2967_n432), 
	.A(n432));
   DLY4X1 FE_PHC2966_plain_text_222_ (.Y(FE_PHN2966_plain_text_222_), 
	.A(FE_PHN1137_plain_text_222_));
   DLY3X1 FE_PHC2965_plain_text_83_ (.Y(FE_PHN2965_plain_text_83_), 
	.A(FE_PHN1146_plain_text_83_));
   DLY3X1 FE_PHC2964_plain_text_148_ (.Y(FE_PHN2964_plain_text_148_), 
	.A(FE_PHN1134_plain_text_148_));
   DLY4X1 FE_PHC2963_n408 (.Y(FE_PHN2963_n408), 
	.A(n408));
   DLY3X1 FE_PHC2962_n469 (.Y(FE_PHN2962_n469), 
	.A(n469));
   DLY4X1 FE_PHC2961_plain_text_45_ (.Y(FE_PHN2961_plain_text_45_), 
	.A(plain_text[45]));
   DLY4X1 FE_PHC2960_plain_text_111_ (.Y(FE_PHN2960_plain_text_111_), 
	.A(plain_text[111]));
   DLY4X1 FE_PHC2959_plain_text_63_ (.Y(FE_PHN2959_plain_text_63_), 
	.A(plain_text[63]));
   DLY3X1 FE_PHC2958_plain_text_88_ (.Y(FE_PHN2958_plain_text_88_), 
	.A(FE_PHN1143_plain_text_88_));
   DLY3X1 FE_PHC2957_plain_text_105_ (.Y(FE_PHN2957_plain_text_105_), 
	.A(plain_text[105]));
   DLY3X1 FE_PHC2953_plain_text_236_ (.Y(FE_PHN2953_plain_text_236_), 
	.A(FE_PHN1339_plain_text_236_));
   DLY3X1 FE_PHC2952_plain_text_97_ (.Y(FE_PHN2952_plain_text_97_), 
	.A(FE_PHN1116_plain_text_97_));
   DLY3X1 FE_PHC2950_plain_text_44_ (.Y(FE_PHN2950_plain_text_44_), 
	.A(FE_PHN1332_plain_text_44_));
   DLY4X1 FE_PHC2949_plain_text_108_ (.Y(FE_PHN2949_plain_text_108_), 
	.A(plain_text[108]));
   DLY4X1 FE_PHC2948_plain_text_119_ (.Y(FE_PHN2948_plain_text_119_), 
	.A(FE_PHN1104_plain_text_119_));
   DLY4X1 FE_PHC2945_plain_text_113_ (.Y(FE_PHN2945_plain_text_113_), 
	.A(FE_PHN1115_plain_text_113_));
   DLY4X1 FE_PHC2944_plain_text_76_ (.Y(FE_PHN2944_plain_text_76_), 
	.A(plain_text[76]));
   DLY3X1 FE_PHC2943_plain_text_151_ (.Y(FE_PHN2943_plain_text_151_), 
	.A(FE_PHN1106_plain_text_151_));
   DLY4X1 FE_PHC2942_plain_text_100_ (.Y(FE_PHN2942_plain_text_100_), 
	.A(FE_PHN1113_plain_text_100_));
   DLY4X1 FE_PHC2940_n510 (.Y(FE_PHN2940_n510), 
	.A(n510));
   DLY4X1 FE_PHC2939_n511 (.Y(FE_PHN2939_n511), 
	.A(n511));
   DLY4X1 FE_PHC2938_n514 (.Y(FE_PHN2938_n514), 
	.A(n514));
   DLY4X1 FE_PHC2937_n512 (.Y(FE_PHN2937_n512), 
	.A(n512));
   DLY4X1 FE_PHC2934_n513 (.Y(FE_PHN2934_n513), 
	.A(n513));
   DLY4X1 FE_PHC2933_plain_text_188_ (.Y(FE_PHN2933_plain_text_188_), 
	.A(plain_text[188]));
   DLY4X1 FE_PHC2932_plain_text_34_ (.Y(FE_PHN2932_plain_text_34_), 
	.A(FE_PHN1316_plain_text_34_));
   DLY4X1 FE_PHC2931_n451 (.Y(FE_PHN2931_n451), 
	.A(n451));
   DLY4X1 FE_PHC2929_plain_text_51_ (.Y(FE_PHN2929_plain_text_51_), 
	.A(FE_PHN1068_plain_text_51_));
   DLY4X1 FE_PHC2928_n457 (.Y(FE_PHN2928_n457), 
	.A(n457));
   DLY4X1 FE_PHC2926_plain_text_53_ (.Y(FE_PHN2926_plain_text_53_), 
	.A(FE_PHN1042_plain_text_53_));
   DLY4X1 FE_PHC2925_plain_text_39_ (.Y(FE_PHN2925_plain_text_39_), 
	.A(FE_PHN1047_plain_text_39_));
   DLY4X1 FE_PHC2924_n509 (.Y(FE_PHN2924_n509), 
	.A(n509));
   DLY2X1 FE_PHC2923_Din_12_ (.Y(plain_key_out[12]), 
	.A(FE_PHN2923_Din_12_));
   DLY2X1 FE_PHC2922_Din_21_ (.Y(plain_key_out[21]), 
	.A(FE_PHN2922_Din_21_));
   DLY4X1 FE_PHC2921_Din_23_ (.Y(plain_key_out[23]), 
	.A(FE_PHN2921_Din_23_));
   DLY3X1 FE_PHC2920_Din_55_ (.Y(plain_key_out[55]), 
	.A(FE_PHN2920_Din_55_));
   DLY3X1 FE_PHC2889_n575 (.Y(FE_PHN2889_n575), 
	.A(n575));
   DLY4X1 FE_PHC2888_plain_text_4_ (.Y(FE_PHN2888_plain_text_4_), 
	.A(FE_PHN888_plain_text_4_));
   DLY3X1 FE_PHC2887_plain_text_155_ (.Y(FE_PHN2887_plain_text_155_), 
	.A(plain_text[155]));
   DLY3X1 FE_PHC2886_n593 (.Y(FE_PHN2886_n593), 
	.A(n593));
   DLY4X1 FE_PHC2885_plain_text_15_ (.Y(FE_PHN2885_plain_text_15_), 
	.A(FE_PHN884_plain_text_15_));
   DLY3X1 FE_PHC2884_plain_text_40_ (.Y(FE_PHN2884_plain_text_40_), 
	.A(FE_PHN1370_plain_text_40_));
   DLY3X1 FE_PHC2883_n626 (.Y(FE_PHN2883_n626), 
	.A(n626));
   DLY4X1 FE_PHC2882_plain_text_77_ (.Y(FE_PHN2882_plain_text_77_), 
	.A(FE_PHN883_plain_text_77_));
   DLY4X1 FE_PHC2881_n688 (.Y(FE_PHN2881_n688), 
	.A(n688));
   DLY4X1 FE_PHC2880_plain_text_16_ (.Y(FE_PHN2880_plain_text_16_), 
	.A(FE_PHN1166_plain_text_16_));
   DLY4X1 FE_PHC2879_n516 (.Y(FE_PHN2879_n516), 
	.A(n516));
   DLY3X1 FE_PHC2878_plain_text_43_ (.Y(FE_PHN2878_plain_text_43_), 
	.A(plain_text[43]));
   DLY3X1 FE_PHC2877_plain_text_134_ (.Y(FE_PHN2877_plain_text_134_), 
	.A(FE_PHN1156_plain_text_134_));
   DLY4X1 FE_PHC2876_plain_text_13_ (.Y(FE_PHN2876_plain_text_13_), 
	.A(FE_PHN874_plain_text_13_));
   DLY4X1 FE_PHC2875_plain_text_36_ (.Y(FE_PHN2875_plain_text_36_), 
	.A(FE_PHN1158_plain_text_36_));
   DLY4X1 FE_PHC2874_plain_text_26_ (.Y(FE_PHN2874_plain_text_26_), 
	.A(FE_PHN875_plain_text_26_));
   DLY4X1 FE_PHC2873_n554 (.Y(FE_PHN2873_n554), 
	.A(n554));
   DLY4X1 FE_PHC2872_n680 (.Y(FE_PHN2872_n680), 
	.A(n680));
   DLY4X1 FE_PHC2871_plain_text_19_ (.Y(FE_PHN2871_plain_text_19_), 
	.A(FE_PHN1150_plain_text_19_));
   DLY3X1 FE_PHC2870_plain_text_239_ (.Y(FE_PHN2870_plain_text_239_), 
	.A(plain_text[239]));
   DLY4X1 FE_PHC2869_n551 (.Y(FE_PHN2869_n551), 
	.A(n551));
   DLY4X1 FE_PHC2868_plain_text_140_ (.Y(FE_PHN2868_plain_text_140_), 
	.A(FE_PHN870_plain_text_140_));
   DLY4X1 FE_PHC2867_plain_text_50_ (.Y(FE_PHN2867_plain_text_50_), 
	.A(FE_PHN1338_plain_text_50_));
   DLY3X1 FE_PHC2866_n669 (.Y(FE_PHN2866_n669), 
	.A(n669));
   DLY4X1 FE_PHC2865_plain_text_62_ (.Y(FE_PHN2865_plain_text_62_), 
	.A(FE_PHN1129_plain_text_62_));
   DLY4X1 FE_PHC2864_n756 (.Y(FE_PHN2864_n756), 
	.A(n756));
   DLY4X1 FE_PHC2863_plain_text_130_ (.Y(FE_PHN2863_plain_text_130_), 
	.A(plain_text[130]));
   DLY4X1 FE_PHC2862_plain_text_143_ (.Y(FE_PHN2862_plain_text_143_), 
	.A(FE_PHN1094_plain_text_143_));
   DLY4X1 FE_PHC2861_plain_text_64_ (.Y(FE_PHN2861_plain_text_64_), 
	.A(FE_PHN1317_plain_text_64_));
   DLY4X1 FE_PHC2860_plain_text_20_ (.Y(FE_PHN2860_plain_text_20_), 
	.A(FE_PHN837_plain_text_20_));
   DLY4X1 FE_PHC2859_n651 (.Y(FE_PHN2859_n651), 
	.A(n651));
   DLY4X1 FE_PHC2858_n636 (.Y(FE_PHN2858_n636), 
	.A(n636));
   DLY4X1 FE_PHC2857_plain_text_197_ (.Y(FE_PHN2857_plain_text_197_), 
	.A(FE_PHN829_plain_text_197_));
   DLY4X1 FE_PHC2854_n739 (.Y(FE_PHN2854_n739), 
	.A(n739));
   DLY4X1 FE_PHC2853_n674 (.Y(FE_PHN2853_n674), 
	.A(n674));
   DLY4X1 FE_PHC2852_n561 (.Y(FE_PHN2852_n561), 
	.A(n561));
   DLY4X1 FE_PHC2851_n711 (.Y(FE_PHN2851_n711), 
	.A(n711));
   BUFXL FE_PHC2822_plain_text_125_ (.Y(FE_PHN2822_plain_text_125_), 
	.A(plain_text[125]));
   DLY2X1 FE_PHC2819_Din_127_ (.Y(plain_key_out[127]), 
	.A(FE_PHN2819_Din_127_));
   DLY2X1 FE_PHC2818_Din_126_ (.Y(plain_key_out[126]), 
	.A(FE_PHN2818_Din_126_));
   DLY2X1 FE_PHC2817_Din_31_ (.Y(plain_key_out[31]), 
	.A(FE_PHN2817_Din_31_));
   DLY4X1 FE_PHC2815_n426 (.Y(FE_PHN2815_n426), 
	.A(n426));
   DLY2X1 FE_PHC2804_pbv1 (.Y(FE_PHN2804_pbv1), 
	.A(pbv1));
   DLY4X1 FE_PHC2801_pf0 (.Y(FE_PHN2801_pf0), 
	.A(pf0));
   DLY4X1 FE_PHC2800_pbv0 (.Y(FE_PHN2800_pbv0), 
	.A(pbv0));
   DLY4X1 FE_PHC2796_n385 (.Y(FE_PHN2796_n385), 
	.A(n385));
   DLY4X1 FE_PHC2794_n474 (.Y(FE_PHN2794_n474), 
	.A(FE_PHN5046_n474));
   DLY4X1 FE_PHC2037_plain_text_124_ (.Y(FE_PHN2037_plain_text_124_), 
	.A(plain_text[124]));
   DLY4X1 FE_PHC2035_plain_text_235_ (.Y(FE_PHN2035_plain_text_235_), 
	.A(FE_PHN3607_plain_text_235_));
   DLY4X1 FE_PHC2034_plain_text_154_ (.Y(FE_PHN2034_plain_text_154_), 
	.A(plain_text[154]));
   DLY4X1 FE_PHC2033_plain_text_238_ (.Y(FE_PHN2033_plain_text_238_), 
	.A(plain_text[238]));
   DLY4X1 FE_PHC2032_plain_text_226_ (.Y(FE_PHN2032_plain_text_226_), 
	.A(plain_text[226]));
   DLY4X1 FE_PHC2031_plain_text_232_ (.Y(FE_PHN2031_plain_text_232_), 
	.A(plain_text[232]));
   DLY4X1 FE_PHC2030_plain_text_219_ (.Y(FE_PHN2030_plain_text_219_), 
	.A(plain_text[219]));
   DLY4X1 FE_PHC2029_plain_text_153_ (.Y(FE_PHN2029_plain_text_153_), 
	.A(FE_PHN5239_plain_text_153_));
   DLY4X1 FE_PHC2028_plain_text_172_ (.Y(FE_PHN2028_plain_text_172_), 
	.A(FE_PHN3597_plain_text_172_));
   DLY4X1 FE_PHC2027_plain_text_184_ (.Y(FE_PHN2027_plain_text_184_), 
	.A(plain_text[184]));
   DLY4X1 FE_PHC2026_plain_text_209_ (.Y(FE_PHN2026_plain_text_209_), 
	.A(plain_text[209]));
   DLY4X1 FE_PHC2025_plain_text_144_ (.Y(FE_PHN2025_plain_text_144_), 
	.A(plain_text[144]));
   DLY4X1 FE_PHC2024_plain_text_165_ (.Y(FE_PHN2024_plain_text_165_), 
	.A(plain_text[165]));
   DLY4X1 FE_PHC2023_plain_text_185_ (.Y(FE_PHN2023_plain_text_185_), 
	.A(FE_PHN5255_plain_text_185_));
   DLY4X1 FE_PHC2022_plain_text_38_ (.Y(FE_PHN2022_plain_text_38_), 
	.A(plain_text[38]));
   DLY4X1 FE_PHC2021_plain_text_229_ (.Y(FE_PHN2021_plain_text_229_), 
	.A(plain_text[229]));
   DLY4X1 FE_PHC2020_plain_text_242_ (.Y(FE_PHN2020_plain_text_242_), 
	.A(plain_text[242]));
   DLY4X1 FE_PHC2019_plain_text_160_ (.Y(FE_PHN2019_plain_text_160_), 
	.A(plain_text[160]));
   DLY4X1 FE_PHC2018_plain_text_204_ (.Y(FE_PHN2018_plain_text_204_), 
	.A(plain_text[204]));
   DLY4X1 FE_PHC2017_plain_text_41_ (.Y(FE_PHN2017_plain_text_41_), 
	.A(plain_text[41]));
   DLY4X1 FE_PHC2016_plain_text_35_ (.Y(FE_PHN2016_plain_text_35_), 
	.A(plain_text[35]));
   DLY4X1 FE_PHC2015_plain_text_67_ (.Y(FE_PHN2015_plain_text_67_), 
	.A(plain_text[67]));
   DLY4X1 FE_PHC2014_plain_text_195_ (.Y(FE_PHN2014_plain_text_195_), 
	.A(plain_text[195]));
   DLY4X1 FE_PHC2013_plain_text_135_ (.Y(FE_PHN2013_plain_text_135_), 
	.A(plain_text[135]));
   DLY4X1 FE_PHC2012_plain_text_233_ (.Y(FE_PHN2012_plain_text_233_), 
	.A(plain_text[233]));
   DLY4X1 FE_PHC2011_plain_text_199_ (.Y(FE_PHN2011_plain_text_199_), 
	.A(plain_text[199]));
   DLY4X1 FE_PHC2010_plain_text_245_ (.Y(FE_PHN2010_plain_text_245_), 
	.A(plain_text[245]));
   DLY4X1 FE_PHC1999_Din_112_ (.Y(plain_key_out[112]), 
	.A(FE_PHN1999_Din_112_));
   DLY4X1 FE_PHC1996_Din_4_ (.Y(plain_key_out[4]), 
	.A(FE_PHN1996_Din_4_));
   DLY4X1 FE_PHC1995_Din_118_ (.Y(plain_key_out[118]), 
	.A(FE_PHN1995_Din_118_));
   DLY4X1 FE_PHC1994_Din_113_ (.Y(plain_key_out[113]), 
	.A(FE_PHN1994_Din_113_));
   DLY4X1 FE_PHC1993_Din_19_ (.Y(plain_key_out[19]), 
	.A(FE_PHN1993_Din_19_));
   DLY4X1 FE_PHC1990_Din_119_ (.Y(plain_key_out[119]), 
	.A(FE_PHN1990_Din_119_));
   DLY4X1 FE_PHC1988_Din_11_ (.Y(plain_key_out[11]), 
	.A(FE_PHN1988_Din_11_));
   DLY4X1 FE_PHC1987_Din_17_ (.Y(plain_key_out[17]), 
	.A(FE_PHN1987_Din_17_));
   DLY4X1 FE_PHC1986_Din_111_ (.Y(plain_key_out[111]), 
	.A(FE_PHN1986_Din_111_));
   DLY4X1 FE_PHC1985_Din_115_ (.Y(plain_key_out[115]), 
	.A(FE_PHN1985_Din_115_));
   DLY4X1 FE_PHC1984_Din_110_ (.Y(plain_key_out[110]), 
	.A(FE_PHN1984_Din_110_));
   DLY4X1 FE_PHC1983_Din_13_ (.Y(plain_key_out[13]), 
	.A(FE_PHN1983_Din_13_));
   DLY4X1 FE_PHC1982_Din_20_ (.Y(plain_key_out[20]), 
	.A(FE_PHN1982_Din_20_));
   DLY4X1 FE_PHC1981_Din_105_ (.Y(plain_key_out[105]), 
	.A(FE_PHN1981_Din_105_));
   DLY4X1 FE_PHC1980_Din_15_ (.Y(plain_key_out[15]), 
	.A(FE_PHN1980_Din_15_));
   DLY4X1 FE_PHC1979_Din_18_ (.Y(plain_key_out[18]), 
	.A(FE_PHN1979_Din_18_));
   DLY4X1 FE_PHC1978_Din_51_ (.Y(plain_key_out[51]), 
	.A(FE_PHN1978_Din_51_));
   DLY4X1 FE_PHC1977_Din_54_ (.Y(plain_key_out[54]), 
	.A(FE_PHN1977_Din_54_));
   DLY4X1 FE_PHC1976_Din_16_ (.Y(plain_key_out[16]), 
	.A(FE_PHN1976_Din_16_));
   DLY4X1 FE_PHC1975_Din_85_ (.Y(plain_key_out[85]), 
	.A(FE_PHN1975_Din_85_));
   DLY4X1 FE_PHC1973_Din_116_ (.Y(plain_key_out[116]), 
	.A(FE_PHN1973_Din_116_));
   DLY4X1 FE_PHC1971_Din_100_ (.Y(plain_key_out[100]), 
	.A(FE_PHN1971_Din_100_));
   DLY4X1 FE_PHC1970_Din_53_ (.Y(plain_key_out[53]), 
	.A(FE_PHN1970_Din_53_));
   DLY4X1 FE_PHC1968_Din_83_ (.Y(plain_key_out[83]), 
	.A(FE_PHN1968_Din_83_));
   DLY4X1 FE_PHC1967_Din_107_ (.Y(plain_key_out[107]), 
	.A(FE_PHN1967_Din_107_));
   DLY4X1 FE_PHC1966_Din_87_ (.Y(plain_key_out[87]), 
	.A(FE_PHN1966_Din_87_));
   DLY4X1 FE_PHC1964_Din_101_ (.Y(plain_key_out[101]), 
	.A(FE_PHN1964_Din_101_));
   DLY4X1 FE_PHC1963_Din_86_ (.Y(plain_key_out[86]), 
	.A(FE_PHN1963_Din_86_));
   DLY4X1 FE_PHC1961_Din_69_ (.Y(plain_key_out[69]), 
	.A(FE_PHN1961_Din_69_));
   DLY4X1 FE_PHC1960_Din_52_ (.Y(plain_key_out[52]), 
	.A(FE_PHN1960_Din_52_));
   DLY4X1 FE_PHC1956_Din_84_ (.Y(plain_key_out[84]), 
	.A(FE_PHN1956_Din_84_));
   DLY4X1 FE_PHC1955_Din_108_ (.Y(plain_key_out[108]), 
	.A(FE_PHN1955_Din_108_));
   DLY4X1 FE_PHC1954_Din_10_ (.Y(plain_key_out[10]), 
	.A(FE_PHN1954_Din_10_));
   DLY4X1 FE_PHC1953_Din_77_ (.Y(plain_key_out[77]), 
	.A(FE_PHN1953_Din_77_));
   DLY4X1 FE_PHC1952_Din_70_ (.Y(plain_key_out[70]), 
	.A(FE_PHN1952_Din_70_));
   DLY4X1 FE_PHC1951_Din_102_ (.Y(plain_key_out[102]), 
	.A(FE_PHN1951_Din_102_));
   DLY4X1 FE_PHC1950_Din_117_ (.Y(plain_key_out[117]), 
	.A(FE_PHN1950_Din_117_));
   DLY4X1 FE_PHC1949_n615 (.Y(FE_PHN1949_n615), 
	.A(n615));
   DLY4X1 FE_PHC1948_Din_109_ (.Y(plain_key_out[109]), 
	.A(FE_PHN1948_Din_109_));
   DLY4X1 FE_PHC1947_n591 (.Y(FE_PHN1947_n591), 
	.A(n591));
   DLY4X1 FE_PHC1946_n517 (.Y(FE_PHN1946_n517), 
	.A(n517));
   DLY4X1 FE_PHC1945_Din_46_ (.Y(plain_key_out[46]), 
	.A(FE_PHN1945_Din_46_));
   DLY4X1 FE_PHC1944_n691 (.Y(FE_PHN1944_n691), 
	.A(n691));
   DLY4X1 FE_PHC1943_Din_78_ (.Y(plain_key_out[78]), 
	.A(FE_PHN1943_Din_78_));
   DLY4X1 FE_PHC1942_Din_37_ (.Y(plain_key_out[37]), 
	.A(FE_PHN1942_Din_37_));
   DLY4X1 FE_PHC1941_Din_45_ (.Y(plain_key_out[45]), 
	.A(FE_PHN1941_Din_45_));
   DLY4X1 FE_PHC1940_Din_43_ (.Y(plain_key_out[43]), 
	.A(FE_PHN1940_Din_43_));
   DLY4X1 FE_PHC1939_n687 (.Y(FE_PHN1939_n687), 
	.A(n687));
   DLY4X1 FE_PHC1938_n528 (.Y(FE_PHN1938_n528), 
	.A(n528));
   DLY4X1 FE_PHC1937_Din_97_ (.Y(plain_key_out[97]), 
	.A(FE_PHN1937_Din_97_));
   DLY4X1 FE_PHC1936_n619 (.Y(FE_PHN1936_n619), 
	.A(n619));
   DLY4X1 FE_PHC1935_n387 (.Y(FE_PHN1935_n387), 
	.A(n387));
   DLY4X1 FE_PHC1934_n660 (.Y(FE_PHN1934_n660), 
	.A(n660));
   DLY4X1 FE_PHC1933_n523 (.Y(FE_PHN1933_n523), 
	.A(n523));
   DLY4X1 FE_PHC1932_n526 (.Y(FE_PHN1932_n526), 
	.A(n526));
   DLY4X1 FE_PHC1931_n555 (.Y(FE_PHN1931_n555), 
	.A(n555));
   DLY4X1 FE_PHC1929_n635 (.Y(FE_PHN1929_n635), 
	.A(n635));
   DLY4X1 FE_PHC1928_n613 (.Y(FE_PHN1928_n613), 
	.A(n613));
   DLY4X1 FE_PHC1927_n678 (.Y(FE_PHN1927_n678), 
	.A(n678));
   DLY4X1 FE_PHC1926_n634 (.Y(FE_PHN1926_n634), 
	.A(n634));
   DLY4X1 FE_PHC1925_Din_103_ (.Y(plain_key_out[103]), 
	.A(FE_PHN1925_Din_103_));
   DLY4X1 FE_PHC1924_n560 (.Y(FE_PHN1924_n560), 
	.A(n560));
   DLY4X1 FE_PHC1923_n618 (.Y(FE_PHN1923_n618), 
	.A(n618));
   DLY4X1 FE_PHC1922_n559 (.Y(FE_PHN1922_n559), 
	.A(n559));
   DLY4X1 FE_PHC1921_n755 (.Y(FE_PHN1921_n755), 
	.A(n755));
   DLY4X1 FE_PHC1920_n583 (.Y(FE_PHN1920_n583), 
	.A(n583));
   DLY4X1 FE_PHC1919_n556 (.Y(FE_PHN1919_n556), 
	.A(n556));
   DLY4X1 FE_PHC1918_n649 (.Y(FE_PHN1918_n649), 
	.A(n649));
   DLY4X1 FE_PHC1916_Din_99_ (.Y(plain_key_out[99]), 
	.A(FE_PHN1916_Din_99_));
   DLY4X1 FE_PHC1915_n573 (.Y(FE_PHN1915_n573), 
	.A(n573));
   DLY4X1 FE_PHC1914_n653 (.Y(FE_PHN1914_n653), 
	.A(n653));
   DLY4X1 FE_PHC1913_Din_75_ (.Y(plain_key_out[75]), 
	.A(FE_PHN1913_Din_75_));
   DLY4X1 FE_PHC1912_n527 (.Y(FE_PHN1912_n527), 
	.A(n527));
   DLY4X1 FE_PHC1911_n735 (.Y(FE_PHN1911_n735), 
	.A(n735));
   DLY4X1 FE_PHC1910_Din_104_ (.Y(plain_key_out[104]), 
	.A(FE_PHN1910_Din_104_));
   DLY4X1 FE_PHC1909_n592 (.Y(FE_PHN1909_n592), 
	.A(n592));
   DLY4X1 FE_PHC1908_Din_82_ (.Y(plain_key_out[82]), 
	.A(FE_PHN1908_Din_82_));
   DLY4X1 FE_PHC1907_Din_76_ (.Y(plain_key_out[76]), 
	.A(FE_PHN1907_Din_76_));
   DLY4X1 FE_PHC1906_n315 (.Y(FE_PHN1906_n315), 
	.A(n315));
   DLY4X1 FE_PHC1904_n283 (.Y(FE_PHN1904_n283), 
	.A(n283));
   DLY4X1 FE_PHC1903_n518 (.Y(FE_PHN1903_n518), 
	.A(n518));
   DLY4X1 FE_PHC1902_n552 (.Y(FE_PHN1902_n552), 
	.A(n552));
   DLY4X1 FE_PHC1901_n281 (.Y(FE_PHN1901_n281), 
	.A(n281));
   DLY4X1 FE_PHC1900_n529 (.Y(FE_PHN1900_n529), 
	.A(n529));
   DLY4X1 FE_PHC1898_n734 (.Y(FE_PHN1898_n734), 
	.A(n734));
   DLY4X1 FE_PHC1897_n291 (.Y(FE_PHN1897_n291), 
	.A(n291));
   DLY4X1 FE_PHC1896_Din_96_ (.Y(plain_key_out[96]), 
	.A(FE_PHN1896_Din_96_));
   DLY4X1 FE_PHC1895_n692 (.Y(FE_PHN1895_n692), 
	.A(n692));
   DLY4X1 FE_PHC1890_n549 (.Y(FE_PHN1890_n549), 
	.A(n549));
   DLY4X1 FE_PHC1886_n524 (.Y(FE_PHN1886_n524), 
	.A(n524));
   DLY4X1 FE_PHC1875_n581 (.Y(FE_PHN1875_n581), 
	.A(n581));
   DLY4X1 FE_PHC1865_n679 (.Y(FE_PHN1865_n679), 
	.A(n679));
   DLY4X1 FE_PHC1845_n553 (.Y(FE_PHN1845_n553), 
	.A(n553));
   DLY4X1 FE_PHC1842_n616 (.Y(FE_PHN1842_n616), 
	.A(n616));
   DLY4X1 FE_PHC1838_plain_text_248_ (.Y(FE_PHN1838_plain_text_248_), 
	.A(plain_text[248]));
   DLY4X1 FE_PHC1836_n550 (.Y(FE_PHN1836_n550), 
	.A(n550));
   DLY4X1 FE_PHC1825_n498 (.Y(FE_PHN1825_n498), 
	.A(n498));
   DLY4X1 FE_PHC1815_n580 (.Y(FE_PHN1815_n580), 
	.A(n580));
   DLY4X1 FE_PHC1753_n574 (.Y(FE_PHN1753_n574), 
	.A(n574));
   DLY4X1 FE_PHC1741_n677 (.Y(FE_PHN1741_n677), 
	.A(n677));
   DLY4X1 FE_PHC1704_n676 (.Y(FE_PHN1704_n676), 
	.A(n676));
   DLY4X1 FE_PHC1465_n747 (.Y(FE_PHN1465_n747), 
	.A(n747));
   DLY4X1 FE_PHC1462_plain_text_1_ (.Y(FE_PHN1462_plain_text_1_), 
	.A(FE_PHN5170_plain_text_1_));
   DLY4X1 FE_PHC1461_plain_text_0_ (.Y(FE_PHN1461_plain_text_0_), 
	.A(plain_text[0]));
   DLY4X1 FE_PHC1460_plain_text_2_ (.Y(FE_PHN1460_plain_text_2_), 
	.A(FE_PHN3181_plain_text_2_));
   DLY4X1 FE_PHC1459_Din_120_ (.Y(plain_key_out[120]), 
	.A(FE_PHN1459_Din_120_));
   DLY4X1 FE_PHC1453_plain_text_5_ (.Y(FE_PHN1453_plain_text_5_), 
	.A(plain_text[5]));
   DLY4X1 FE_PHC1452_plain_text_123_ (.Y(FE_PHN1452_plain_text_123_), 
	.A(FE_PHN3176_plain_text_123_));
   DLY4X1 FE_PHC1451_plain_text_14_ (.Y(FE_PHN1451_plain_text_14_), 
	.A(plain_text[14]));
   DLY4X1 FE_PHC1450_plain_text_6_ (.Y(FE_PHN1450_plain_text_6_), 
	.A(FE_PHN3175_plain_text_6_));
   DLY4X1 FE_PHC1448_plain_text_7_ (.Y(FE_PHN1448_plain_text_7_), 
	.A(plain_text[7]));
   DLY4X1 FE_PHC1447_plain_text_214_ (.Y(FE_PHN1447_plain_text_214_), 
	.A(plain_text[214]));
   DLY4X1 FE_PHC1443_plain_text_182_ (.Y(FE_PHN1443_plain_text_182_), 
	.A(plain_text[182]));
   DLY4X1 FE_PHC1440_plain_text_132_ (.Y(FE_PHN1440_plain_text_132_), 
	.A(plain_text[132]));
   DLY4X1 FE_PHC1439_plain_text_183_ (.Y(FE_PHN1439_plain_text_183_), 
	.A(plain_text[183]));
   DLY4X1 FE_PHC1438_plain_text_122_ (.Y(FE_PHN1438_plain_text_122_), 
	.A(FE_PHN3167_plain_text_122_));
   DLY4X1 FE_PHC1437_n443 (.Y(FE_PHN1437_n443), 
	.A(n443));
   DLY4X1 FE_PHC1436_plain_text_126_ (.Y(FE_PHN1436_plain_text_126_), 
	.A(plain_text[126]));
   DLY4X1 FE_PHC1435_n386 (.Y(FE_PHN1435_n386), 
	.A(n386));
   DLY4X1 FE_PHC1433_plain_text_246_ (.Y(FE_PHN1433_plain_text_246_), 
	.A(plain_text[246]));
   DLY4X1 FE_PHC1432_plain_text_215_ (.Y(FE_PHN1432_plain_text_215_), 
	.A(plain_text[215]));
   DLY4X1 FE_PHC1431_n475 (.Y(FE_PHN1431_n475), 
	.A(FE_PHN5048_n475));
   DLY4X1 FE_PHC1430_plain_text_179_ (.Y(FE_PHN1430_plain_text_179_), 
	.A(FE_PHN3166_plain_text_179_));
   DLY4X1 FE_PHC1428_plain_text_69_ (.Y(FE_PHN1428_plain_text_69_), 
	.A(plain_text[69]));
   DLY4X1 FE_PHC1427_plain_text_147_ (.Y(FE_PHN1427_plain_text_147_), 
	.A(FE_PHN3390_plain_text_147_));
   DLY4X1 FE_PHC1426_plain_text_25_ (.Y(FE_PHN1426_plain_text_25_), 
	.A(plain_text[25]));
   DLY4X1 FE_PHC1424_plain_text_12_ (.Y(FE_PHN1424_plain_text_12_), 
	.A(plain_text[12]));
   DLY4X1 FE_PHC1423_n272 (.Y(FE_PHN1423_n272), 
	.A(n272));
   DLY4X1 FE_PHC1420_plain_text_189_ (.Y(FE_PHN1420_plain_text_189_), 
	.A(plain_text[189]));
   DLY4X1 FE_PHC1418_plain_text_205_ (.Y(FE_PHN1418_plain_text_205_), 
	.A(plain_text[205]));
   DLY4X1 FE_PHC1417_plain_text_187_ (.Y(FE_PHN1417_plain_text_187_), 
	.A(plain_text[187]));
   DLY4X1 FE_PHC1411_plain_text_171_ (.Y(FE_PHN1411_plain_text_171_), 
	.A(FE_PHN3156_plain_text_171_));
   DLY4X1 FE_PHC1410_plain_text_28_ (.Y(FE_PHN1410_plain_text_28_), 
	.A(plain_text[28]));
   DLY4X1 FE_PHC1409_plain_text_210_ (.Y(FE_PHN1409_plain_text_210_), 
	.A(plain_text[210]));
   DLY4X1 FE_PHC1407_n486 (.Y(FE_PHN1407_n486), 
	.A(n486));
   DLY4X1 FE_PHC1403_plain_text_174_ (.Y(FE_PHN1403_plain_text_174_), 
	.A(plain_text[174]));
   DLY4X1 FE_PHC1400_plain_text_240_ (.Y(FE_PHN1400_plain_text_240_), 
	.A(plain_text[240]));
   DLY4X1 FE_PHC1399_plain_text_138_ (.Y(FE_PHN1399_plain_text_138_), 
	.A(plain_text[138]));
   DLY4X1 FE_PHC1398_plain_text_228_ (.Y(FE_PHN1398_plain_text_228_), 
	.A(FE_PHN3162_plain_text_228_));
   DLY4X1 FE_PHC1396_plain_text_145_ (.Y(FE_PHN1396_plain_text_145_), 
	.A(plain_text[145]));
   DLY4X1 FE_PHC1390_plain_text_178_ (.Y(FE_PHN1390_plain_text_178_), 
	.A(plain_text[178]));
   DLY4X1 FE_PHC1389_plain_text_218_ (.Y(FE_PHN1389_plain_text_218_), 
	.A(plain_text[218]));
   DLY4X1 FE_PHC1387_plain_text_139_ (.Y(FE_PHN1387_plain_text_139_), 
	.A(plain_text[139]));
   DLY4X1 FE_PHC1386_plain_text_200_ (.Y(FE_PHN1386_plain_text_200_), 
	.A(plain_text[200]));
   DLY4X1 FE_PHC1385_plain_text_177_ (.Y(FE_PHN1385_plain_text_177_), 
	.A(plain_text[177]));
   DLY4X1 FE_PHC1384_plain_text_58_ (.Y(FE_PHN1384_plain_text_58_), 
	.A(FE_PHN3063_plain_text_58_));
   DLY4X1 FE_PHC1383_plain_text_18_ (.Y(FE_PHN1383_plain_text_18_), 
	.A(plain_text[18]));
   DLY4X1 FE_PHC1382_plain_text_48_ (.Y(FE_PHN1382_plain_text_48_), 
	.A(FE_PHN3151_plain_text_48_));
   DLY4X1 FE_PHC1381_plain_text_216_ (.Y(FE_PHN1381_plain_text_216_), 
	.A(plain_text[216]));
   DLY4X1 FE_PHC1379_plain_text_163_ (.Y(FE_PHN1379_plain_text_163_), 
	.A(plain_text[163]));
   DLY4X1 FE_PHC1378_plain_text_196_ (.Y(FE_PHN1378_plain_text_196_), 
	.A(plain_text[196]));
   DLY4X1 FE_PHC1377_plain_text_30_ (.Y(FE_PHN1377_plain_text_30_), 
	.A(plain_text[30]));
   DLY4X1 FE_PHC1376_plain_text_194_ (.Y(FE_PHN1376_plain_text_194_), 
	.A(plain_text[194]));
   DLY4X1 FE_PHC1374_plain_text_231_ (.Y(FE_PHN1374_plain_text_231_), 
	.A(FE_PHN3157_plain_text_231_));
   DLY4X1 FE_PHC1373_plain_text_202_ (.Y(FE_PHN1373_plain_text_202_), 
	.A(plain_text[202]));
   DLY4X1 FE_PHC1372_plain_text_206_ (.Y(FE_PHN1372_plain_text_206_), 
	.A(plain_text[206]));
   DLY4X1 FE_PHC1371_plain_text_169_ (.Y(FE_PHN1371_plain_text_169_), 
	.A(plain_text[169]));
   DLY4X1 FE_PHC1370_plain_text_40_ (.Y(FE_PHN1370_plain_text_40_), 
	.A(plain_text[40]));
   DLY4X1 FE_PHC1369_plain_text_65_ (.Y(FE_PHN1369_plain_text_65_), 
	.A(FE_PHN3146_plain_text_65_));
   DLY4X1 FE_PHC1368_plain_text_224_ (.Y(FE_PHN1368_plain_text_224_), 
	.A(plain_text[224]));
   DLY4X1 FE_PHC1366_plain_text_114_ (.Y(FE_PHN1366_plain_text_114_), 
	.A(plain_text[114]));
   DLY4X1 FE_PHC1365_plain_text_170_ (.Y(FE_PHN1365_plain_text_170_), 
	.A(FE_PHN3133_plain_text_170_));
   DLY4X1 FE_PHC1364_plain_text_136_ (.Y(FE_PHN1364_plain_text_136_), 
	.A(plain_text[136]));
   DLY4X1 FE_PHC1363_plain_text_175_ (.Y(FE_PHN1363_plain_text_175_), 
	.A(plain_text[175]));
   DLY4X1 FE_PHC1362_plain_text_72_ (.Y(FE_PHN1362_plain_text_72_), 
	.A(plain_text[72]));
   DLY4X1 FE_PHC1361_plain_text_243_ (.Y(FE_PHN1361_plain_text_243_), 
	.A(plain_text[243]));
   DLY4X1 FE_PHC1359_plain_text_42_ (.Y(FE_PHN1359_plain_text_42_), 
	.A(FE_PHN3400_plain_text_42_));
   DLY4X1 FE_PHC1358_plain_text_198_ (.Y(FE_PHN1358_plain_text_198_), 
	.A(FE_PHN3139_plain_text_198_));
   DLY4X1 FE_PHC1357_n423 (.Y(FE_PHN1357_n423), 
	.A(n423));
   DLY4X1 FE_PHC1356_n456 (.Y(FE_PHN1356_n456), 
	.A(n456));
   DLY4X1 FE_PHC1355_plain_text_32_ (.Y(FE_PHN1355_plain_text_32_), 
	.A(FE_PHN3404_plain_text_32_));
   DLY4X1 FE_PHC1354_plain_text_98_ (.Y(FE_PHN1354_plain_text_98_), 
	.A(plain_text[98]));
   DLY4X1 FE_PHC1352_plain_text_79_ (.Y(FE_PHN1352_plain_text_79_), 
	.A(plain_text[79]));
   DLY4X1 FE_PHC1351_plain_text_213_ (.Y(FE_PHN1351_plain_text_213_), 
	.A(plain_text[213]));
   DLY4X1 FE_PHC1350_plain_text_176_ (.Y(FE_PHN1350_plain_text_176_), 
	.A(plain_text[176]));
   DLY4X1 FE_PHC1349_plain_text_71_ (.Y(FE_PHN1349_plain_text_71_), 
	.A(FE_PHN3002_plain_text_71_));
   DLY4X1 FE_PHC1348_plain_text_80_ (.Y(FE_PHN1348_plain_text_80_), 
	.A(plain_text[80]));
   DLY4X1 FE_PHC1347_plain_text_129_ (.Y(FE_PHN1347_plain_text_129_), 
	.A(plain_text[129]));
   DLY4X1 FE_PHC1346_plain_text_230_ (.Y(FE_PHN1346_plain_text_230_), 
	.A(plain_text[230]));
   DLY4X1 FE_PHC1344_plain_text_73_ (.Y(FE_PHN1344_plain_text_73_), 
	.A(FE_PHN3048_plain_text_73_));
   DLY4X1 FE_PHC1343_plain_text_81_ (.Y(FE_PHN1343_plain_text_81_), 
	.A(FE_PHN3128_plain_text_81_));
   DLY4X1 FE_PHC1342_plain_text_74_ (.Y(FE_PHN1342_plain_text_74_), 
	.A(FE_PHN2985_plain_text_74_));
   DLY4X1 FE_PHC1341_plain_text_142_ (.Y(FE_PHN1341_plain_text_142_), 
	.A(plain_text[142]));
   DLY4X1 FE_PHC1340_n721 (.Y(FE_PHN1340_n721), 
	.A(n721));
   DLY4X1 FE_PHC1339_plain_text_236_ (.Y(FE_PHN1339_plain_text_236_), 
	.A(plain_text[236]));
   DLY4X1 FE_PHC1338_plain_text_50_ (.Y(FE_PHN1338_plain_text_50_), 
	.A(plain_text[50]));
   DLY4X1 FE_PHC1337_plain_text_128_ (.Y(FE_PHN1337_plain_text_128_), 
	.A(plain_text[128]));
   DLY4X1 FE_PHC1336_plain_text_239_ (.Y(FE_PHN1336_plain_text_239_), 
	.A(FE_PHN2870_plain_text_239_));
   DLY4X1 FE_PHC1334_plain_text_47_ (.Y(FE_PHN1334_plain_text_47_), 
	.A(FE_PHN3110_plain_text_47_));
   DLY4X1 FE_PHC1332_plain_text_44_ (.Y(FE_PHN1332_plain_text_44_), 
	.A(plain_text[44]));
   DLY4X1 FE_PHC1331_plain_text_244_ (.Y(FE_PHN1331_plain_text_244_), 
	.A(plain_text[244]));
   DLY4X1 FE_PHC1330_n425 (.Y(FE_PHN1330_n425), 
	.A(n425));
   DLY4X1 FE_PHC1329_plain_text_201_ (.Y(FE_PHN1329_plain_text_201_), 
	.A(plain_text[201]));
   DLY4X1 FE_PHC1328_plain_text_106_ (.Y(FE_PHN1328_plain_text_106_), 
	.A(FE_PHN5236_plain_text_106_));
   DLY4X1 FE_PHC1327_plain_text_141_ (.Y(FE_PHN1327_plain_text_141_), 
	.A(FE_PHN3126_plain_text_141_));
   DLY4X1 FE_PHC1325_plain_text_137_ (.Y(FE_PHN1325_plain_text_137_), 
	.A(FE_PHN3114_plain_text_137_));
   DLY4X1 FE_PHC1320_plain_text_68_ (.Y(FE_PHN1320_plain_text_68_), 
	.A(FE_PHN3125_plain_text_68_));
   DLY4X1 FE_PHC1319_n508 (.Y(FE_PHN1319_n508), 
	.A(n508));
   DLY4X1 FE_PHC1317_plain_text_64_ (.Y(FE_PHN1317_plain_text_64_), 
	.A(plain_text[64]));
   DLY4X1 FE_PHC1316_plain_text_34_ (.Y(FE_PHN1316_plain_text_34_), 
	.A(plain_text[34]));
   DLY4X1 FE_PHC1309_Din_5_ (.Y(plain_key_out[5]), 
	.A(FE_PHN1309_Din_5_));
   DLY4X1 FE_PHC1308_Din_2_ (.Y(plain_key_out[2]), 
	.A(FE_PHN1308_Din_2_));
   DLY4X1 FE_PHC1307_Din_1_ (.Y(plain_key_out[1]), 
	.A(FE_PHN1307_Din_1_));
   DLY4X1 FE_PHC1306_Din_38_ (.Y(plain_key_out[38]), 
	.A(FE_PHN1306_Din_38_));
   DLY4X1 FE_PHC1305_Din_3_ (.Y(plain_key_out[3]), 
	.A(FE_PHN1305_Din_3_));
   DLY4X1 FE_PHC1304_Din_0_ (.Y(plain_key_out[0]), 
	.A(FE_PHN1304_Din_0_));
   DLY4X1 FE_PHC1303_Din_36_ (.Y(plain_key_out[36]), 
	.A(FE_PHN1303_Din_36_));
   DLY4X1 FE_PHC1302_Din_7_ (.Y(plain_key_out[7]), 
	.A(FE_PHN1302_Din_7_));
   DLY4X1 FE_PHC1301_Din_67_ (.Y(plain_key_out[67]), 
	.A(FE_PHN1301_Din_67_));
   DLY4X1 FE_PHC1300_Din_68_ (.Y(plain_key_out[68]), 
	.A(FE_PHN1300_Din_68_));
   DLY4X1 FE_PHC1298_Din_35_ (.Y(plain_key_out[35]), 
	.A(FE_PHN1298_Din_35_));
   DLY4X1 FE_PHC1297_Din_71_ (.Y(plain_key_out[71]), 
	.A(FE_PHN1297_Din_71_));
   DLY4X1 FE_PHC1296_Din_66_ (.Y(plain_key_out[66]), 
	.A(FE_PHN1296_Din_66_));
   DLY4X1 FE_PHC1295_Din_6_ (.Y(plain_key_out[6]), 
	.A(FE_PHN1295_Din_6_));
   DLY4X1 FE_PHC1294_Din_44_ (.Y(plain_key_out[44]), 
	.A(FE_PHN1294_Din_44_));
   DLY4X1 FE_PHC1293_Din_64_ (.Y(plain_key_out[64]), 
	.A(FE_PHN1293_Din_64_));
   DLY4X1 FE_PHC1292_Din_48_ (.Y(plain_key_out[48]), 
	.A(FE_PHN1292_Din_48_));
   DLY4X1 FE_PHC1291_Din_80_ (.Y(plain_key_out[80]), 
	.A(FE_PHN1291_Din_80_));
   DLY4X1 FE_PHC1290_Din_73_ (.Y(plain_key_out[73]), 
	.A(FE_PHN1290_Din_73_));
   DLY4X1 FE_PHC1287_Din_74_ (.Y(plain_key_out[74]), 
	.A(FE_PHN1287_Din_74_));
   DLY4X1 FE_PHC1286_Din_50_ (.Y(plain_key_out[50]), 
	.A(FE_PHN1286_Din_50_));
   DLY4X1 FE_PHC1285_Din_40_ (.Y(plain_key_out[40]), 
	.A(FE_PHN1285_Din_40_));
   DLY4X1 FE_PHC1283_Din_65_ (.Y(plain_key_out[65]), 
	.A(FE_PHN1283_Din_65_));
   DLY4X1 FE_PHC1282_Din_106_ (.Y(plain_key_out[106]), 
	.A(FE_PHN1282_Din_106_));
   DLY4X1 FE_PHC1281_Din_81_ (.Y(plain_key_out[81]), 
	.A(FE_PHN1281_Din_81_));
   DLY4X1 FE_PHC1280_Din_42_ (.Y(plain_key_out[42]), 
	.A(FE_PHN1280_Din_42_));
   DLY4X1 FE_PHC1279_Din_22_ (.Y(plain_key_out[22]), 
	.A(FE_PHN1279_Din_22_));
   DLY4X1 FE_PHC1278_Din_114_ (.Y(plain_key_out[114]), 
	.A(FE_PHN1278_Din_114_));
   DLY4X1 FE_PHC1277_Din_39_ (.Y(plain_key_out[39]), 
	.A(FE_PHN1277_Din_39_));
   DLY4X1 FE_PHC1276_Din_79_ (.Y(plain_key_out[79]), 
	.A(FE_PHN1276_Din_79_));
   DLY4X1 FE_PHC1275_Din_49_ (.Y(plain_key_out[49]), 
	.A(FE_PHN1275_Din_49_));
   DLY4X1 FE_PHC1274_Din_98_ (.Y(plain_key_out[98]), 
	.A(FE_PHN1274_Din_98_));
   DLY4X1 FE_PHC1273_Din_41_ (.Y(plain_key_out[41]), 
	.A(FE_PHN1273_Din_41_));
   DLY4X1 FE_PHC1272_Din_9_ (.Y(plain_key_out[9]), 
	.A(FE_PHN1272_Din_9_));
   DLY4X1 FE_PHC1271_Din_34_ (.Y(plain_key_out[34]), 
	.A(FE_PHN1271_Din_34_));
   DLY4X1 FE_PHC1270_Din_32_ (.Y(plain_key_out[32]), 
	.A(FE_PHN1270_Din_32_));
   DLY4X1 FE_PHC1269_Din_14_ (.Y(plain_key_out[14]), 
	.A(FE_PHN1269_Din_14_));
   DLY4X1 FE_PHC1268_Din_8_ (.Y(plain_key_out[8]), 
	.A(FE_PHN1268_Din_8_));
   DLY4X1 FE_PHC1267_Din_47_ (.Y(plain_key_out[47]), 
	.A(FE_PHN1267_Din_47_));
   DLY4X1 FE_PHC1266_Din_72_ (.Y(plain_key_out[72]), 
	.A(FE_PHN1266_Din_72_));
   DLY4X1 FE_PHC1260_Din_33_ (.Y(plain_key_out[33]), 
	.A(FE_PHN1260_Din_33_));
   DLY4X1 FE_PHC1250_plain_text_251_ (.Y(FE_PHN1250_plain_text_251_), 
	.A(FE_PHN3088_plain_text_251_));
   DLY4X1 FE_PHC1248_plain_text_254_ (.Y(FE_PHN1248_plain_text_254_), 
	.A(plain_text[254]));
   DLY4X1 FE_PHC1243_n812 (.Y(FE_PHN1243_n812), 
	.A(n812));
   DLY4X1 FE_PHC1242_plain_text_250_ (.Y(FE_PHN1242_plain_text_250_), 
	.A(plain_text[250]));
   DLY4X1 FE_PHC1240_plain_text_252_ (.Y(FE_PHN1240_plain_text_252_), 
	.A(plain_text[252]));
   DLY4X1 FE_PHC1228_plain_text_253_ (.Y(FE_PHN1228_plain_text_253_), 
	.A(plain_text[253]));
   DLY4X1 FE_PHC1218_plain_text_249_ (.Y(FE_PHN1218_plain_text_249_), 
	.A(FE_PHN3082_plain_text_249_));
   DLY4X1 FE_PHC1217_Din_121_ (.Y(plain_key_out[121]), 
	.A(FE_PHN1217_Din_121_));
   DLY4X1 FE_PHC1216_Din_27_ (.Y(plain_key_out[27]), 
	.A(FE_PHN1216_Din_27_));
   DLY4X1 FE_PHC1215_Din_28_ (.Y(plain_key_out[28]), 
	.A(FE_PHN1215_Din_28_));
   DLY4X1 FE_PHC1214_Din_29_ (.Y(plain_key_out[29]), 
	.A(FE_PHN1214_Din_29_));
   DLY4X1 FE_PHC1213_Din_123_ (.Y(plain_key_out[123]), 
	.A(FE_PHN1213_Din_123_));
   DLY4X1 FE_PHC1212_n659 (.Y(FE_PHN1212_n659), 
	.A(n659));
   DLY4X1 FE_PHC1210_plain_text_3_ (.Y(FE_PHN1210_plain_text_3_), 
	.A(FE_PHN3074_plain_text_3_));
   DLY4X1 FE_PHC1209_plain_text_157_ (.Y(FE_PHN1209_plain_text_157_), 
	.A(plain_text[157]));
   DLY4X1 FE_PHC1208_plain_text_133_ (.Y(FE_PHN1208_plain_text_133_), 
	.A(plain_text[133]));
   DLY4X1 FE_PHC1207_plain_text_118_ (.Y(FE_PHN1207_plain_text_118_), 
	.A(plain_text[118]));
   DLY4X1 FE_PHC1206_plain_text_116_ (.Y(FE_PHN1206_plain_text_116_), 
	.A(plain_text[116]));
   DLY4X1 FE_PHC1205_plain_text_24_ (.Y(FE_PHN1205_plain_text_24_), 
	.A(plain_text[24]));
   DLY4X1 FE_PHC1204_plain_text_59_ (.Y(FE_PHN1204_plain_text_59_), 
	.A(plain_text[59]));
   DLY4X1 FE_PHC1203_n546 (.Y(FE_PHN1203_n546), 
	.A(n546));
   DLY4X1 FE_PHC1202_plain_text_17_ (.Y(FE_PHN1202_plain_text_17_), 
	.A(plain_text[17]));
   DLY4X1 FE_PHC1201_plain_text_8_ (.Y(FE_PHN1201_plain_text_8_), 
	.A(plain_text[8]));
   DLY4X1 FE_PHC1200_plain_text_109_ (.Y(FE_PHN1200_plain_text_109_), 
	.A(plain_text[109]));
   DLY4X1 FE_PHC1199_plain_text_127_ (.Y(FE_PHN1199_plain_text_127_), 
	.A(plain_text[127]));
   DLY4X1 FE_PHC1198_n625 (.Y(FE_PHN1198_n625), 
	.A(n625));
   DLY4X1 FE_PHC1196_plain_text_54_ (.Y(FE_PHN1196_plain_text_54_), 
	.A(FE_PHN3141_plain_text_54_));
   DLY4X1 FE_PHC1195_plain_text_162_ (.Y(FE_PHN1195_plain_text_162_), 
	.A(plain_text[162]));
   DLY4X1 FE_PHC1194_plain_text_152_ (.Y(FE_PHN1194_plain_text_152_), 
	.A(plain_text[152]));
   DLY4X1 FE_PHC1193_plain_text_101_ (.Y(FE_PHN1193_plain_text_101_), 
	.A(plain_text[101]));
   DLY4X1 FE_PHC1192_plain_text_22_ (.Y(FE_PHN1192_plain_text_22_), 
	.A(plain_text[22]));
   DLY4X1 FE_PHC1191_plain_text_150_ (.Y(FE_PHN1191_plain_text_150_), 
	.A(plain_text[150]));
   DLY4X1 FE_PHC1190_plain_text_146_ (.Y(FE_PHN1190_plain_text_146_), 
	.A(plain_text[146]));
   DLY4X1 FE_PHC1189_plain_text_70_ (.Y(FE_PHN1189_plain_text_70_), 
	.A(plain_text[70]));
   DLY4X1 FE_PHC1188_plain_text_121_ (.Y(FE_PHN1188_plain_text_121_), 
	.A(FE_PHN5154_plain_text_121_));
   DLY4X1 FE_PHC1187_plain_text_61_ (.Y(FE_PHN1187_plain_text_61_), 
	.A(FE_PHN3011_plain_text_61_));
   DLY4X1 FE_PHC1186_n609 (.Y(FE_PHN1186_n609), 
	.A(n609));
   DLY4X1 FE_PHC1185_plain_text_186_ (.Y(FE_PHN1185_plain_text_186_), 
	.A(plain_text[186]));
   DLY4X1 FE_PHC1184_plain_text_92_ (.Y(FE_PHN1184_plain_text_92_), 
	.A(plain_text[92]));
   DLY4X1 FE_PHC1183_plain_text_223_ (.Y(FE_PHN1183_plain_text_223_), 
	.A(plain_text[223]));
   DLY4X1 FE_PHC1182_plain_text_91_ (.Y(FE_PHN1182_plain_text_91_), 
	.A(plain_text[91]));
   DLY4X1 FE_PHC1181_plain_text_78_ (.Y(FE_PHN1181_plain_text_78_), 
	.A(FE_PHN5243_plain_text_78_));
   DLY4X1 FE_PHC1180_plain_text_203_ (.Y(FE_PHN1180_plain_text_203_), 
	.A(FE_PHN3350_plain_text_203_));
   DLY4X1 FE_PHC1179_plain_text_208_ (.Y(FE_PHN1179_plain_text_208_), 
	.A(plain_text[208]));
   DLY4X1 FE_PHC1178_plain_text_85_ (.Y(FE_PHN1178_plain_text_85_), 
	.A(plain_text[85]));
   DLY4X1 FE_PHC1177_plain_text_112_ (.Y(FE_PHN1177_plain_text_112_), 
	.A(plain_text[112]));
   DLY4X1 FE_PHC1176_plain_text_60_ (.Y(FE_PHN1176_plain_text_60_), 
	.A(FE_PHN3098_plain_text_60_));
   DLY4X1 FE_PHC1175_plain_text_99_ (.Y(FE_PHN1175_plain_text_99_), 
	.A(plain_text[99]));
   DLY4X1 FE_PHC1174_plain_text_159_ (.Y(FE_PHN1174_plain_text_159_), 
	.A(plain_text[159]));
   DLY4X1 FE_PHC1173_plain_text_117_ (.Y(FE_PHN1173_plain_text_117_), 
	.A(plain_text[117]));
   DLY4X1 FE_PHC1171_plain_text_86_ (.Y(FE_PHN1171_plain_text_86_), 
	.A(plain_text[86]));
   DLY4X1 FE_PHC1170_plain_text_11_ (.Y(FE_PHN1170_plain_text_11_), 
	.A(FE_PHN3163_plain_text_11_));
   DLY4X1 FE_PHC1169_plain_text_181_ (.Y(FE_PHN1169_plain_text_181_), 
	.A(FE_PHN2989_plain_text_181_));
   DLY4X1 FE_PHC1168_plain_text_173_ (.Y(FE_PHN1168_plain_text_173_), 
	.A(FE_PHN2988_plain_text_173_));
   DLY4X1 FE_PHC1167_plain_text_93_ (.Y(FE_PHN1167_plain_text_93_), 
	.A(FE_PHN3051_plain_text_93_));
   DLY4X1 FE_PHC1166_plain_text_16_ (.Y(FE_PHN1166_plain_text_16_), 
	.A(plain_text[16]));
   DLY4X1 FE_PHC1165_plain_text_190_ (.Y(FE_PHN1165_plain_text_190_), 
	.A(plain_text[190]));
   DLY4X1 FE_PHC1163_plain_text_168_ (.Y(FE_PHN1163_plain_text_168_), 
	.A(FE_PHN3354_plain_text_168_));
   DLY4X1 FE_PHC1162_plain_text_149_ (.Y(FE_PHN1162_plain_text_149_), 
	.A(plain_text[149]));
   DLY4X1 FE_PHC1161_plain_text_193_ (.Y(FE_PHN1161_plain_text_193_), 
	.A(plain_text[193]));
   DLY4X1 FE_PHC1160_plain_text_156_ (.Y(FE_PHN1160_plain_text_156_), 
	.A(FE_PHN3007_plain_text_156_));
   DLY4X1 FE_PHC1159_plain_text_37_ (.Y(FE_PHN1159_plain_text_37_), 
	.A(plain_text[37]));
   DLY4X1 FE_PHC1158_plain_text_36_ (.Y(FE_PHN1158_plain_text_36_), 
	.A(plain_text[36]));
   DLY4X1 FE_PHC1157_plain_text_29_ (.Y(FE_PHN1157_plain_text_29_), 
	.A(plain_text[29]));
   DLY4X1 FE_PHC1156_plain_text_134_ (.Y(FE_PHN1156_plain_text_134_), 
	.A(plain_text[134]));
   DLY4X1 FE_PHC1155_plain_text_9_ (.Y(FE_PHN1155_plain_text_9_), 
	.A(plain_text[9]));
   DLY4X1 FE_PHC1154_n459 (.Y(FE_PHN1154_n459), 
	.A(n459));
   DLY4X1 FE_PHC1153_plain_text_95_ (.Y(FE_PHN1153_plain_text_95_), 
	.A(FE_PHN3041_plain_text_95_));
   DLY4X1 FE_PHC1152_plain_text_158_ (.Y(FE_PHN1152_plain_text_158_), 
	.A(FE_PHN2984_plain_text_158_));
   DLY4X1 FE_PHC1151_plain_text_107_ (.Y(FE_PHN1151_plain_text_107_), 
	.A(plain_text[107]));
   DLY4X1 FE_PHC1150_plain_text_19_ (.Y(FE_PHN1150_plain_text_19_), 
	.A(plain_text[19]));
   DLY4X1 FE_PHC1149_plain_text_45_ (.Y(FE_PHN1149_plain_text_45_), 
	.A(FE_PHN2961_plain_text_45_));
   DLY4X1 FE_PHC1148_plain_text_120_ (.Y(FE_PHN1148_plain_text_120_), 
	.A(FE_PHN3032_plain_text_120_));
   DLY4X1 FE_PHC1147_plain_text_241_ (.Y(FE_PHN1147_plain_text_241_), 
	.A(FE_PHN3337_plain_text_241_));
   DLY4X1 FE_PHC1146_plain_text_83_ (.Y(FE_PHN1146_plain_text_83_), 
	.A(plain_text[83]));
   DLY4X1 FE_PHC1145_plain_text_115_ (.Y(FE_PHN1145_plain_text_115_), 
	.A(FE_PHN3019_plain_text_115_));
   DLY4X1 FE_PHC1144_plain_text_131_ (.Y(FE_PHN1144_plain_text_131_), 
	.A(plain_text[131]));
   DLY4X1 FE_PHC1143_plain_text_88_ (.Y(FE_PHN1143_plain_text_88_), 
	.A(plain_text[88]));
   DLY4X1 FE_PHC1142_plain_text_89_ (.Y(FE_PHN1142_plain_text_89_), 
	.A(FE_PHN3009_plain_text_89_));
   DLY4X1 FE_PHC1141_plain_text_90_ (.Y(FE_PHN1141_plain_text_90_), 
	.A(plain_text[90]));
   DLY4X1 FE_PHC1140_n710 (.Y(FE_PHN1140_n710), 
	.A(n710));
   DLY4X1 FE_PHC1139_plain_text_234_ (.Y(FE_PHN1139_plain_text_234_), 
	.A(plain_text[234]));
   DLY4X1 FE_PHC1138_plain_text_55_ (.Y(FE_PHN1138_plain_text_55_), 
	.A(FE_PHN3320_plain_text_55_));
   DLY4X1 FE_PHC1137_plain_text_222_ (.Y(FE_PHN1137_plain_text_222_), 
	.A(plain_text[222]));
   DLY4X1 FE_PHC1136_n395 (.Y(FE_PHN1136_n395), 
	.A(n395));
   DLY4X1 FE_PHC1135_plain_text_102_ (.Y(FE_PHN1135_plain_text_102_), 
	.A(plain_text[102]));
   DLY4X1 FE_PHC1134_plain_text_148_ (.Y(FE_PHN1134_plain_text_148_), 
	.A(plain_text[148]));
   DLY4X1 FE_PHC1133_plain_text_21_ (.Y(FE_PHN1133_plain_text_21_), 
	.A(FE_PHN3280_plain_text_21_));
   DLY4X1 FE_PHC1132_plain_text_207_ (.Y(FE_PHN1132_plain_text_207_), 
	.A(FE_PHN3023_plain_text_207_));
   DLY4X1 FE_PHC1131_plain_text_63_ (.Y(FE_PHN1131_plain_text_63_), 
	.A(FE_PHN2959_plain_text_63_));
   DLY4X1 FE_PHC1130_plain_text_221_ (.Y(FE_PHN1130_plain_text_221_), 
	.A(plain_text[221]));
   DLY4X1 FE_PHC1129_plain_text_62_ (.Y(FE_PHN1129_plain_text_62_), 
	.A(plain_text[62]));
   DLY4X1 FE_PHC1128_n434 (.Y(FE_PHN1128_n434), 
	.A(n434));
   DLY4X1 FE_PHC1127_plain_text_161_ (.Y(FE_PHN1127_plain_text_161_), 
	.A(FE_PHN3298_plain_text_161_));
   DLY4X1 FE_PHC1126_plain_text_31_ (.Y(FE_PHN1126_plain_text_31_), 
	.A(FE_PHN3299_plain_text_31_));
   DLY4X1 FE_PHC1125_plain_text_23_ (.Y(FE_PHN1125_plain_text_23_), 
	.A(FE_PHN3318_plain_text_23_));
   DLY4X1 FE_PHC1124_plain_text_130_ (.Y(FE_PHN1124_plain_text_130_), 
	.A(FE_PHN2863_plain_text_130_));
   DLY4X1 FE_PHC1123_plain_text_110_ (.Y(FE_PHN1123_plain_text_110_), 
	.A(plain_text[110]));
   DLY4X1 FE_PHC1122_plain_text_56_ (.Y(FE_PHN1122_plain_text_56_), 
	.A(FE_PHN3135_plain_text_56_));
   DLY4X1 FE_PHC1121_n725 (.Y(FE_PHN1121_n725), 
	.A(n725));
   DLY4X1 FE_PHC1120_plain_text_108_ (.Y(FE_PHN1120_plain_text_108_), 
	.A(FE_PHN2949_plain_text_108_));
   DLY4X1 FE_PHC1119_plain_text_84_ (.Y(FE_PHN1119_plain_text_84_), 
	.A(FE_PHN3006_plain_text_84_));
   DLY4X1 FE_PHC1118_plain_text_211_ (.Y(FE_PHN1118_plain_text_211_), 
	.A(plain_text[211]));
   DLY4X1 FE_PHC1117_plain_text_225_ (.Y(FE_PHN1117_plain_text_225_), 
	.A(plain_text[225]));
   DLY4X1 FE_PHC1116_plain_text_97_ (.Y(FE_PHN1116_plain_text_97_), 
	.A(plain_text[97]));
   DLY4X1 FE_PHC1115_plain_text_113_ (.Y(FE_PHN1115_plain_text_113_), 
	.A(plain_text[113]));
   DLY4X1 FE_PHC1114_plain_text_66_ (.Y(FE_PHN1114_plain_text_66_), 
	.A(FE_PHN3005_plain_text_66_));
   DLY4X1 FE_PHC1113_plain_text_100_ (.Y(FE_PHN1113_plain_text_100_), 
	.A(plain_text[100]));
   DLY4X1 FE_PHC1112_plain_text_104_ (.Y(FE_PHN1112_plain_text_104_), 
	.A(FE_PHN2979_plain_text_104_));
   DLY4X1 FE_PHC1111_plain_text_57_ (.Y(FE_PHN1111_plain_text_57_), 
	.A(FE_PHN2999_plain_text_57_));
   DLY4X1 FE_PHC1110_plain_text_103_ (.Y(FE_PHN1110_plain_text_103_), 
	.A(FE_PHN3033_plain_text_103_));
   DLY4X1 FE_PHC1109_plain_text_96_ (.Y(FE_PHN1109_plain_text_96_), 
	.A(plain_text[96]));
   DLY4X1 FE_PHC1108_plain_text_192_ (.Y(FE_PHN1108_plain_text_192_), 
	.A(FE_PHN3287_plain_text_192_));
   DLY4X1 FE_PHC1106_plain_text_151_ (.Y(FE_PHN1106_plain_text_151_), 
	.A(plain_text[151]));
   DLY4X1 FE_PHC1105_plain_text_220_ (.Y(FE_PHN1105_plain_text_220_), 
	.A(FE_PHN2968_plain_text_220_));
   DLY4X1 FE_PHC1104_plain_text_119_ (.Y(FE_PHN1104_plain_text_119_), 
	.A(plain_text[119]));
   DLY4X1 FE_PHC1103_plain_text_76_ (.Y(FE_PHN1103_plain_text_76_), 
	.A(FE_PHN2944_plain_text_76_));
   DLY4X1 FE_PHC1102_plain_text_164_ (.Y(FE_PHN1102_plain_text_164_), 
	.A(FE_PHN2976_plain_text_164_));
   DLY4X1 FE_PHC1101_plain_text_87_ (.Y(FE_PHN1101_plain_text_87_), 
	.A(FE_PHN2972_plain_text_87_));
   DLY4X1 FE_PHC1099_plain_text_217_ (.Y(FE_PHN1099_plain_text_217_), 
	.A(FE_PHN3093_plain_text_217_));
   DLY4X1 FE_PHC1097_plain_text_82_ (.Y(FE_PHN1097_plain_text_82_), 
	.A(FE_PHN3001_plain_text_82_));
   DLY4X1 FE_PHC1095_plain_text_94_ (.Y(FE_PHN1095_plain_text_94_), 
	.A(FE_PHN2980_plain_text_94_));
   DLY4X1 FE_PHC1094_plain_text_143_ (.Y(FE_PHN1094_plain_text_143_), 
	.A(plain_text[143]));
   DLY4X1 FE_PHC1091_plain_text_27_ (.Y(FE_PHN1091_plain_text_27_), 
	.A(plain_text[27]));
   DLY4X1 FE_PHC1090_n639 (.Y(FE_PHN1090_n639), 
	.A(n639));
   DLY4X1 FE_PHC1089_plain_text_49_ (.Y(FE_PHN1089_plain_text_49_), 
	.A(FE_PHN3090_plain_text_49_));
   DLY4X1 FE_PHC1082_plain_text_33_ (.Y(FE_PHN1082_plain_text_33_), 
	.A(FE_PHN3379_plain_text_33_));
   DLY4X1 FE_PHC1078_plain_text_105_ (.Y(FE_PHN1078_plain_text_105_), 
	.A(FE_PHN2957_plain_text_105_));
   DLY4X1 FE_PHC1073_plain_text_52_ (.Y(FE_PHN1073_plain_text_52_), 
	.A(FE_PHN3348_plain_text_52_));
   DLY4X1 FE_PHC1072_n668 (.Y(FE_PHN1072_n668), 
	.A(n668));
   DLY4X1 FE_PHC1071_plain_text_111_ (.Y(FE_PHN1071_plain_text_111_), 
	.A(FE_PHN2960_plain_text_111_));
   DLY4X1 FE_PHC1070_n740 (.Y(FE_PHN1070_n740), 
	.A(n740));
   DLY4X1 FE_PHC1069_plain_text_247_ (.Y(FE_PHN1069_plain_text_247_), 
	.A(plain_text[247]));
   DLY4X1 FE_PHC1068_plain_text_51_ (.Y(FE_PHN1068_plain_text_51_), 
	.A(plain_text[51]));
   DLY4X1 FE_PHC1065_plain_text_167_ (.Y(FE_PHN1065_plain_text_167_), 
	.A(plain_text[167]));
   DLY4X1 FE_PHC1061_n644 (.Y(FE_PHN1061_n644), 
	.A(n644));
   DLY4X1 FE_PHC1059_plain_text_188_ (.Y(FE_PHN1059_plain_text_188_), 
	.A(FE_PHN2933_plain_text_188_));
   DLY4X1 FE_PHC1047_plain_text_39_ (.Y(FE_PHN1047_plain_text_39_), 
	.A(plain_text[39]));
   DLY4X1 FE_PHC1042_plain_text_53_ (.Y(FE_PHN1042_plain_text_53_), 
	.A(plain_text[53]));
   DLY4X1 FE_PHC1039_plain_text_166_ (.Y(FE_PHN1039_plain_text_166_), 
	.A(plain_text[166]));
   DLY4X1 FE_PHC911_Din_93_ (.Y(plain_key_out[93]), 
	.A(FE_PHN911_Din_93_));
   DLY4X1 FE_PHC910_Din_24_ (.Y(plain_key_out[24]), 
	.A(FE_PHN910_Din_24_));
   DLY4X1 FE_PHC909_Din_124_ (.Y(plain_key_out[124]), 
	.A(FE_PHN909_Din_124_));
   DLY4X1 FE_PHC908_Din_26_ (.Y(plain_key_out[26]), 
	.A(FE_PHN908_Din_26_));
   DLY4X1 FE_PHC907_Din_25_ (.Y(plain_key_out[25]), 
	.A(FE_PHN907_Din_25_));
   DLY4X1 FE_PHC906_Din_94_ (.Y(plain_key_out[94]), 
	.A(FE_PHN906_Din_94_));
   DLY4X1 FE_PHC904_Din_88_ (.Y(plain_key_out[88]), 
	.A(FE_PHN904_Din_88_));
   DLY4X1 FE_PHC903_Din_56_ (.Y(plain_key_out[56]), 
	.A(FE_PHN903_Din_56_));
   DLY4X1 FE_PHC902_Din_122_ (.Y(plain_key_out[122]), 
	.A(FE_PHN902_Din_122_));
   DLY4X1 FE_PHC901_Din_59_ (.Y(plain_key_out[59]), 
	.A(FE_PHN901_Din_59_));
   DLY4X1 FE_PHC900_Din_91_ (.Y(plain_key_out[91]), 
	.A(FE_PHN900_Din_91_));
   DLY4X1 FE_PHC899_Din_60_ (.Y(plain_key_out[60]), 
	.A(FE_PHN899_Din_60_));
   DLY4X1 FE_PHC898_Din_57_ (.Y(plain_key_out[57]), 
	.A(FE_PHN898_Din_57_));
   DLY4X1 FE_PHC897_Din_90_ (.Y(plain_key_out[90]), 
	.A(FE_PHN897_Din_90_));
   DLY4X1 FE_PHC895_Din_63_ (.Y(plain_key_out[63]), 
	.A(FE_PHN895_Din_63_));
   DLY4X1 FE_PHC894_Din_62_ (.Y(plain_key_out[62]), 
	.A(FE_PHN894_Din_62_));
   DLY4X1 FE_PHC893_Din_58_ (.Y(plain_key_out[58]), 
	.A(FE_PHN893_Din_58_));
   DLY4X1 FE_PHC892_Din_61_ (.Y(plain_key_out[61]), 
	.A(FE_PHN892_Din_61_));
   DLY4X1 FE_PHC891_Din_95_ (.Y(plain_key_out[95]), 
	.A(FE_PHN891_Din_95_));
   DLY4X1 FE_PHC890_Din_89_ (.Y(plain_key_out[89]), 
	.A(FE_PHN890_Din_89_));
   DLY4X1 FE_PHC889_Din_92_ (.Y(plain_key_out[92]), 
	.A(FE_PHN889_Din_92_));
   DLY4X1 FE_PHC888_plain_text_4_ (.Y(FE_PHN888_plain_text_4_), 
	.A(plain_text[4]));
   DLY4X1 FE_PHC886_plain_text_227_ (.Y(FE_PHN886_plain_text_227_), 
	.A(plain_text[227]));
   DLY4X1 FE_PHC884_plain_text_15_ (.Y(FE_PHN884_plain_text_15_), 
	.A(plain_text[15]));
   DLY4X1 FE_PHC883_plain_text_77_ (.Y(FE_PHN883_plain_text_77_), 
	.A(plain_text[77]));
   DLY4X1 FE_PHC882_plain_text_155_ (.Y(FE_PHN882_plain_text_155_), 
	.A(FE_PHN2887_plain_text_155_));
   DLY4X1 FE_PHC880_plain_text_10_ (.Y(FE_PHN880_plain_text_10_), 
	.A(plain_text[10]));
   DLY4X1 FE_PHC875_plain_text_26_ (.Y(FE_PHN875_plain_text_26_), 
	.A(plain_text[26]));
   DLY4X1 FE_PHC874_plain_text_13_ (.Y(FE_PHN874_plain_text_13_), 
	.A(plain_text[13]));
   DLY4X1 FE_PHC870_plain_text_140_ (.Y(FE_PHN870_plain_text_140_), 
	.A(plain_text[140]));
   DLY4X1 FE_PHC864_plain_text_43_ (.Y(FE_PHN864_plain_text_43_), 
	.A(FE_PHN2878_plain_text_43_));
   DLY4X1 FE_PHC861_plain_text_75_ (.Y(FE_PHN861_plain_text_75_), 
	.A(plain_text[75]));
   DLY4X1 FE_PHC860_plain_text_212_ (.Y(FE_PHN860_plain_text_212_), 
	.A(FE_PHN3100_plain_text_212_));
   DLY4X1 FE_PHC837_plain_text_20_ (.Y(FE_PHN837_plain_text_20_), 
	.A(plain_text[20]));
   DLY4X1 FE_PHC835_plain_text_237_ (.Y(FE_PHN835_plain_text_237_), 
	.A(plain_text[237]));
   DLY4X1 FE_PHC830_plain_text_180_ (.Y(FE_PHN830_plain_text_180_), 
	.A(FE_PHN3086_plain_text_180_));
   DLY4X1 FE_PHC829_plain_text_197_ (.Y(FE_PHN829_plain_text_197_), 
	.A(plain_text[197]));
   DLY4X1 FE_PHC828_plain_text_46_ (.Y(FE_PHN828_plain_text_46_), 
	.A(FE_PHN3083_plain_text_46_));
   DLY4X1 FE_PHC824_plain_text_191_ (.Y(FE_PHN824_plain_text_191_), 
	.A(plain_text[191]));
   DLY4X1 FE_PHC823_n718 (.Y(FE_PHN823_n718), 
	.A(n718));
   DLY4X1 FE_PHC749_Din_125_ (.Y(plain_key_out[125]), 
	.A(FE_PHN749_Din_125_));
   DLY4X1 FE_PHC742_Din_30_ (.Y(plain_key_out[30]), 
	.A(FE_PHN742_Din_30_));
   DLY4X1 FE_PHC711_n427 (.Y(FE_PHN711_n427), 
	.A(n427));
   DLY4X1 FE_PHC704_n258 (.Y(FE_PHN704_n258), 
	.A(n258));
   DLY4X1 FE_PHC680_Din_183_ (.Y(plain_key_out[183]), 
	.A(FE_PHN680_Din_183_));
   DLY4X1 FE_PHC679_Din_182_ (.Y(plain_key_out[182]), 
	.A(FE_PHN679_Din_182_));
   DLY4X1 FE_PHC677_Din_158_ (.Y(plain_key_out[158]), 
	.A(FE_PHN677_Din_158_));
   DLY4X1 FE_PHC676_Din_157_ (.Y(plain_key_out[157]), 
	.A(FE_PHN676_Din_157_));
   DLY4X1 FE_PHC675_Din_155_ (.Y(plain_key_out[155]), 
	.A(FE_PHN675_Din_155_));
   DLY4X1 FE_PHC674_Din_147_ (.Y(plain_key_out[147]), 
	.A(FE_PHN674_Din_147_));
   DLY4X1 FE_PHC673_Din_148_ (.Y(plain_key_out[148]), 
	.A(FE_PHN673_Din_148_));
   DLY4X1 FE_PHC672_Din_156_ (.Y(plain_key_out[156]), 
	.A(FE_PHN672_Din_156_));
   DLY4X1 FE_PHC671_Din_149_ (.Y(plain_key_out[149]), 
	.A(FE_PHN671_Din_149_));
   DLY4X1 FE_PHC670_Din_211_ (.Y(plain_key_out[211]), 
	.A(FE_PHN670_Din_211_));
   DLY4X1 FE_PHC669_Din_146_ (.Y(plain_key_out[146]), 
	.A(FE_PHN669_Din_146_));
   DLY4X1 FE_PHC668_Din_186_ (.Y(plain_key_out[186]), 
	.A(FE_PHN668_Din_186_));
   DLY4X1 FE_PHC667_Din_159_ (.Y(plain_key_out[159]), 
	.A(FE_PHN667_Din_159_));
   DLY4X1 FE_PHC666_Din_180_ (.Y(plain_key_out[180]), 
	.A(FE_PHN666_Din_180_));
   DLY4X1 FE_PHC665_Din_188_ (.Y(plain_key_out[188]), 
	.A(FE_PHN665_Din_188_));
   DLY4X1 FE_PHC664_Din_250_ (.Y(plain_key_out[250]), 
	.A(FE_PHN664_Din_250_));
   DLY4X1 FE_PHC663_Din_225_ (.Y(plain_key_out[225]), 
	.A(FE_PHN663_Din_225_));
   DLY4X1 FE_PHC662_Din_208_ (.Y(plain_key_out[208]), 
	.A(FE_PHN662_Din_208_));
   DLY4X1 FE_PHC661_Din_181_ (.Y(plain_key_out[181]), 
	.A(FE_PHN661_Din_181_));
   DLY4X1 FE_PHC660_Din_151_ (.Y(plain_key_out[151]), 
	.A(FE_PHN660_Din_151_));
   DLY4X1 FE_PHC659_Din_247_ (.Y(plain_key_out[247]), 
	.A(FE_PHN659_Din_247_));
   DLY4X1 FE_PHC658_Din_252_ (.Y(plain_key_out[252]), 
	.A(FE_PHN658_Din_252_));
   DLY4X1 FE_PHC657_Din_212_ (.Y(plain_key_out[212]), 
	.A(FE_PHN657_Din_212_));
   DLY4X1 FE_PHC656_Din_150_ (.Y(plain_key_out[150]), 
	.A(FE_PHN656_Din_150_));
   DLY4X1 FE_PHC655_Din_140_ (.Y(plain_key_out[140]), 
	.A(FE_PHN655_Din_140_));
   DLY4X1 FE_PHC654_Din_220_ (.Y(plain_key_out[220]), 
	.A(FE_PHN654_Din_220_));
   DLY4X1 FE_PHC653_Din_227_ (.Y(plain_key_out[227]), 
	.A(FE_PHN653_Din_227_));
   DLY4X1 FE_PHC652_Din_237_ (.Y(plain_key_out[237]), 
	.A(FE_PHN652_Din_237_));
   DLY4X1 FE_PHC651_Din_221_ (.Y(plain_key_out[221]), 
	.A(FE_PHN651_Din_221_));
   DLY4X1 FE_PHC650_Din_249_ (.Y(plain_key_out[249]), 
	.A(FE_PHN650_Din_249_));
   DLY4X1 FE_PHC649_Din_244_ (.Y(plain_key_out[244]), 
	.A(FE_PHN649_Din_244_));
   DLY4X1 FE_PHC648_Din_241_ (.Y(plain_key_out[241]), 
	.A(FE_PHN5230_Din_241_));
   DLY4X1 FE_PHC647_Din_255_ (.Y(plain_key_out[255]), 
	.A(FE_PHN647_Din_255_));
   DLY4X1 FE_PHC645_Din_251_ (.Y(plain_key_out[251]), 
	.A(FE_PHN645_Din_251_));
   DLY4X1 FE_PHC644_Din_166_ (.Y(plain_key_out[166]), 
	.A(FE_PHN644_Din_166_));
   DLY4X1 FE_PHC643_Din_164_ (.Y(plain_key_out[164]), 
	.A(FE_PHN643_Din_164_));
   DLY4X1 FE_PHC642_Din_253_ (.Y(plain_key_out[253]), 
	.A(FE_PHN642_Din_253_));
   DLY4X1 FE_PHC641_Din_191_ (.Y(plain_key_out[191]), 
	.A(FE_PHN641_Din_191_));
   DLY4X1 FE_PHC640_Din_254_ (.Y(plain_key_out[254]), 
	.A(FE_PHN640_Din_254_));
   DLY4X1 FE_PHC639_Din_197_ (.Y(plain_key_out[197]), 
	.A(FE_PHN639_Din_197_));
   DLY4X1 FE_PHC637_Din_167_ (.Y(plain_key_out[167]), 
	.A(FE_PHN637_Din_167_));
   DLY4X1 FE_PHC532_Din_219_ (.Y(plain_key_out[219]), 
	.A(FE_PHN532_Din_219_));
   DLY4X1 FE_PHC531_Din_139_ (.Y(plain_key_out[139]), 
	.A(FE_PHN531_Din_139_));
   DLY4X1 FE_PHC530_Din_154_ (.Y(plain_key_out[154]), 
	.A(FE_PHN530_Din_154_));
   DLY4X1 FE_PHC529_Din_189_ (.Y(plain_key_out[189]), 
	.A(FE_PHN529_Din_189_));
   DLY4X1 FE_PHC527_Din_187_ (.Y(plain_key_out[187]), 
	.A(FE_PHN527_Din_187_));
   DLY4X1 FE_PHC526_Din_210_ (.Y(plain_key_out[210]), 
	.A(FE_PHN526_Din_210_));
   DLY4X1 FE_PHC525_Din_202_ (.Y(plain_key_out[202]), 
	.A(FE_PHN525_Din_202_));
   DLY4X1 FE_PHC524_Din_228_ (.Y(plain_key_out[228]), 
	.A(FE_PHN524_Din_228_));
   DLY4X1 FE_PHC523_Din_160_ (.Y(plain_key_out[160]), 
	.A(FE_PHN523_Din_160_));
   DLY4X1 FE_PHC522_Din_246_ (.Y(plain_key_out[246]), 
	.A(FE_PHN522_Din_246_));
   DLY4X1 FE_PHC521_Din_130_ (.Y(plain_key_out[130]), 
	.A(FE_PHN521_Din_130_));
   DLY4X1 FE_PHC520_Din_226_ (.Y(plain_key_out[226]), 
	.A(FE_PHN520_Din_226_));
   DLY4X1 FE_PHC519_Din_185_ (.Y(plain_key_out[185]), 
	.A(FE_PHN519_Din_185_));
   DLY4X1 FE_PHC518_Din_153_ (.Y(plain_key_out[153]), 
	.A(FE_PHN518_Din_153_));
   DLY4X1 FE_PHC517_Din_236_ (.Y(plain_key_out[236]), 
	.A(FE_PHN517_Din_236_));
   DLY4X1 FE_PHC516_Din_231_ (.Y(plain_key_out[231]), 
	.A(FE_PHN516_Din_231_));
   DLY4X1 FE_PHC515_Din_134_ (.Y(plain_key_out[134]), 
	.A(FE_PHN515_Din_134_));
   DLY4X1 FE_PHC514_Din_218_ (.Y(plain_key_out[218]), 
	.A(FE_PHN514_Din_218_));
   DLY4X1 FE_PHC513_Din_203_ (.Y(plain_key_out[203]), 
	.A(FE_PHN513_Din_203_));
   DLY4X1 FE_PHC512_Din_200_ (.Y(plain_key_out[200]), 
	.A(FE_PHN512_Din_200_));
   DLY4X1 FE_PHC511_Din_141_ (.Y(plain_key_out[141]), 
	.A(FE_PHN511_Din_141_));
   DLY4X1 FE_PHC510_Din_177_ (.Y(plain_key_out[177]), 
	.A(FE_PHN510_Din_177_));
   DLY4X1 FE_PHC509_Din_204_ (.Y(plain_key_out[204]), 
	.A(FE_PHN509_Din_204_));
   DLY4X1 FE_PHC508_Din_195_ (.Y(plain_key_out[195]), 
	.A(FE_PHN508_Din_195_));
   DLY4X1 FE_PHC507_Din_213_ (.Y(plain_key_out[213]), 
	.A(FE_PHN507_Din_213_));
   DLY4X1 FE_PHC506_Din_178_ (.Y(plain_key_out[178]), 
	.A(FE_PHN506_Din_178_));
   DLY4X1 FE_PHC504_Din_179_ (.Y(plain_key_out[179]), 
	.A(FE_PHN504_Din_179_));
   DLY4X1 FE_PHC503_Din_142_ (.Y(plain_key_out[142]), 
	.A(FE_PHN503_Din_142_));
   DLY4X1 FE_PHC502_Din_184_ (.Y(plain_key_out[184]), 
	.A(FE_PHN502_Din_184_));
   DLY4X1 FE_PHC501_Din_222_ (.Y(plain_key_out[222]), 
	.A(FE_PHN501_Din_222_));
   DLY4X1 FE_PHC500_Din_217_ (.Y(plain_key_out[217]), 
	.A(FE_PHN500_Din_217_));
   DLY4X1 FE_PHC499_Din_229_ (.Y(plain_key_out[229]), 
	.A(FE_PHN499_Din_229_));
   DLY4X1 FE_PHC498_Din_233_ (.Y(plain_key_out[233]), 
	.A(FE_PHN498_Din_233_));
   DLY4X1 FE_PHC497_Din_205_ (.Y(plain_key_out[205]), 
	.A(FE_PHN497_Din_205_));
   DLY4X1 FE_PHC496_Din_173_ (.Y(plain_key_out[173]), 
	.A(FE_PHN496_Din_173_));
   DLY4X1 FE_PHC495_Din_162_ (.Y(plain_key_out[162]), 
	.A(FE_PHN495_Din_162_));
   DLY4X1 FE_PHC494_Din_196_ (.Y(plain_key_out[196]), 
	.A(FE_PHN494_Din_196_));
   DLY4X1 FE_PHC493_Din_163_ (.Y(plain_key_out[163]), 
	.A(FE_PHN493_Din_163_));
   DLY4X1 FE_PHC492_Din_224_ (.Y(plain_key_out[224]), 
	.A(FE_PHN492_Din_224_));
   DLY4X1 FE_PHC491_Din_152_ (.Y(plain_key_out[152]), 
	.A(FE_PHN491_Din_152_));
   DLY4X1 FE_PHC490_Din_234_ (.Y(plain_key_out[234]), 
	.A(FE_PHN490_Din_234_));
   DLY4X1 FE_PHC489_Din_199_ (.Y(plain_key_out[199]), 
	.A(FE_PHN489_Din_199_));
   DLY4X1 FE_PHC488_Din_168_ (.Y(plain_key_out[168]), 
	.A(FE_PHN488_Din_168_));
   DLY4X1 FE_PHC487_Din_194_ (.Y(plain_key_out[194]), 
	.A(FE_PHN487_Din_194_));
   DLY4X1 FE_PHC486_Din_243_ (.Y(plain_key_out[243]), 
	.A(FE_PHN486_Din_243_));
   DLY4X1 FE_PHC485_Din_176_ (.Y(plain_key_out[176]), 
	.A(FE_PHN485_Din_176_));
   DLY4X1 FE_PHC484_Din_169_ (.Y(plain_key_out[169]), 
	.A(FE_PHN484_Din_169_));
   DLY4X1 FE_PHC483_Din_230_ (.Y(plain_key_out[230]), 
	.A(FE_PHN483_Din_230_));
   DLY4X1 FE_PHC482_Din_135_ (.Y(plain_key_out[135]), 
	.A(FE_PHN482_Din_135_));
   DLY4X1 FE_PHC481_Din_190_ (.Y(plain_key_out[190]), 
	.A(FE_PHN481_Din_190_));
   DLY4X1 FE_PHC480_Din_239_ (.Y(plain_key_out[239]), 
	.A(FE_PHN480_Din_239_));
   DLY4X1 FE_PHC479_Din_193_ (.Y(plain_key_out[193]), 
	.A(FE_PHN479_Din_193_));
   DLY4X1 FE_PHC478_Din_192_ (.Y(plain_key_out[192]), 
	.A(FE_PHN478_Din_192_));
   DLY4X1 FE_PHC477_Din_235_ (.Y(plain_key_out[235]), 
	.A(FE_PHN477_Din_235_));
   DLY4X1 FE_PHC476_Din_245_ (.Y(plain_key_out[245]), 
	.A(FE_PHN476_Din_245_));
   DLY4X1 FE_PHC475_Din_223_ (.Y(plain_key_out[223]), 
	.A(FE_PHN475_Din_223_));
   DLY4X1 FE_PHC474_Din_242_ (.Y(plain_key_out[242]), 
	.A(FE_PHN474_Din_242_));
   DLY4X1 FE_PHC473_Din_138_ (.Y(plain_key_out[138]), 
	.A(FE_PHN473_Din_138_));
   DLY4X1 FE_PHC472_Din_174_ (.Y(plain_key_out[174]), 
	.A(FE_PHN472_Din_174_));
   DLY4X1 FE_PHC471_Din_145_ (.Y(plain_key_out[145]), 
	.A(FE_PHN471_Din_145_));
   DLY4X1 FE_PHC470_Din_206_ (.Y(plain_key_out[206]), 
	.A(FE_PHN470_Din_206_));
   DLY4X1 FE_PHC469_Din_207_ (.Y(plain_key_out[207]), 
	.A(FE_PHN469_Din_207_));
   DLY4X1 FE_PHC468_Din_171_ (.Y(plain_key_out[171]), 
	.A(FE_PHN468_Din_171_));
   DLY4X1 FE_PHC467_Din_201_ (.Y(plain_key_out[201]), 
	.A(FE_PHN467_Din_201_));
   DLY4X1 FE_PHC466_Din_144_ (.Y(plain_key_out[144]), 
	.A(FE_PHN466_Din_144_));
   DLY4X1 FE_PHC465_Din_165_ (.Y(plain_key_out[165]), 
	.A(FE_PHN465_Din_165_));
   DLY4X1 FE_PHC464_Din_216_ (.Y(plain_key_out[216]), 
	.A(FE_PHN464_Din_216_));
   DLY4X1 FE_PHC463_Din_170_ (.Y(plain_key_out[170]), 
	.A(FE_PHN463_Din_170_));
   DLY4X1 FE_PHC462_Din_128_ (.Y(plain_key_out[128]), 
	.A(FE_PHN462_Din_128_));
   DLY4X1 FE_PHC461_Din_136_ (.Y(plain_key_out[136]), 
	.A(FE_PHN461_Din_136_));
   DLY4X1 FE_PHC460_Din_143_ (.Y(plain_key_out[143]), 
	.A(FE_PHN460_Din_143_));
   DLY4X1 FE_PHC459_Din_238_ (.Y(plain_key_out[238]), 
	.A(FE_PHN459_Din_238_));
   DLY4X1 FE_PHC458_Din_131_ (.Y(plain_key_out[131]), 
	.A(FE_PHN458_Din_131_));
   DLY4X1 FE_PHC457_Din_129_ (.Y(plain_key_out[129]), 
	.A(FE_PHN457_Din_129_));
   DLY4X1 FE_PHC456_Din_232_ (.Y(plain_key_out[232]), 
	.A(FE_PHN456_Din_232_));
   DLY4X1 FE_PHC455_Din_209_ (.Y(plain_key_out[209]), 
	.A(FE_PHN455_Din_209_));
   DLY4X1 FE_PHC454_Din_198_ (.Y(plain_key_out[198]), 
	.A(FE_PHN454_Din_198_));
   DLY4X1 FE_PHC453_Din_240_ (.Y(plain_key_out[240]), 
	.A(FE_PHN453_Din_240_));
   DLY4X1 FE_PHC452_Din_172_ (.Y(plain_key_out[172]), 
	.A(FE_PHN452_Din_172_));
   DLY4X1 FE_PHC451_Din_133_ (.Y(plain_key_out[133]), 
	.A(FE_PHN451_Din_133_));
   DLY4X1 FE_PHC450_Din_161_ (.Y(plain_key_out[161]), 
	.A(FE_PHN450_Din_161_));
   DLY4X1 FE_PHC449_Din_132_ (.Y(plain_key_out[132]), 
	.A(FE_PHN449_Din_132_));
   DLY4X1 FE_PHC448_Din_137_ (.Y(plain_key_out[137]), 
	.A(FE_PHN448_Din_137_));
   DLY4X1 FE_PHC447_Din_175_ (.Y(plain_key_out[175]), 
	.A(FE_PHN447_Din_175_));
   DLY4X1 FE_PHC446_Din_248_ (.Y(plain_key_out[248]), 
	.A(FE_PHN446_Din_248_));
   CLKBUFX2 FE_PHC119_n1 (.Y(FE_PHN119_n1), 
	.A(n1));
   CLKINVX2 FE_OFC75_n1 (.Y(FE_OFN75_n1), 
	.A(FE_OFN67_n1));
   CLKINVX2 FE_OFC74_n1 (.Y(FE_OFN74_n1), 
	.A(FE_OFN67_n1));
   CLKINVX2 FE_OFC73_n1 (.Y(FE_OFN73_n1), 
	.A(FE_OFN67_n1));
   INVX2 FE_OFC72_n1 (.Y(FE_OFN72_n1), 
	.A(FE_OFN67_n1));
   INVX1 FE_OFC71_n1 (.Y(FE_OFN71_n1), 
	.A(FE_OFN67_n1));
   CLKINVX2 FE_OFC70_n1 (.Y(FE_OFN70_n1), 
	.A(FE_OFN67_n1));
   CLKINVX2 FE_OFC69_n1 (.Y(FE_OFN69_n1), 
	.A(FE_OFN67_n1));
   CLKBUFX2 FE_OFC68_n1 (.Y(FE_OFN68_n1), 
	.A(FE_PHN119_n1));
   INVX1 FE_OFC67_n1 (.Y(FE_OFN67_n1), 
	.A(FE_PHN119_n1));
   CLKBUFX3 FE_OFC66_n258 (.Y(FE_OFN66_n258), 
	.A(FE_OFN65_n258));
   CLKBUFX3 FE_OFC65_n258 (.Y(FE_OFN65_n258), 
	.A(FE_OFN64_n258));
   CLKBUFX3 FE_OFC64_n258 (.Y(FE_OFN64_n258), 
	.A(FE_PHN704_n258));
   CLKINVX3 FE_OFC63_n210 (.Y(FE_OFN63_n210), 
	.A(FE_OFN59_n210));
   CLKINVX3 FE_OFC62_n210 (.Y(FE_OFN62_n210), 
	.A(FE_OFN59_n210));
   INVX2 FE_OFC61_n210 (.Y(FE_OFN61_n210), 
	.A(FE_OFN59_n210));
   INVX2 FE_OFC60_n210 (.Y(FE_OFN60_n210), 
	.A(FE_OFN59_n210));
   INVX1 FE_OFC59_n210 (.Y(FE_OFN59_n210), 
	.A(n210));
   CLKBUFX2 FE_OFC52_reset_n (.Y(FE_OFN52_reset_n), 
	.A(FE_OFN42_reset_n));
   DFFRHQX1 plain_text_reg_7_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[7]), 
	.D(FE_PHN3170_n771), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 plain_text_reg_15_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[15]), 
	.D(n770), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_23_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[23]), 
	.D(n769), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_31_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[31]), 
	.D(FE_PHN3317_n768), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_39_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[39]), 
	.D(n767), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_47_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[47]), 
	.D(n766), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_55_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[55]), 
	.D(FE_PHN3254_n765), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_63_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[63]), 
	.D(n764), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_71_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[71]), 
	.D(n763), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_79_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[79]), 
	.D(n762), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_87_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[87]), 
	.D(n761), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_95_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[95]), 
	.D(n760), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_103_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[103]), 
	.D(n759), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_111_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[111]), 
	.D(n758), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_119_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[119]), 
	.D(n757), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_127_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[127]), 
	.D(FE_PHN2864_n756), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_135_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[135]), 
	.D(FE_PHN1921_n755), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_143_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[143]), 
	.D(FE_PHN3127_n754), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_151_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[151]), 
	.D(n753), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_159_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[159]), 
	.D(n752), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_167_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[167]), 
	.D(FE_PHN3120_n751), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_175_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[175]), 
	.D(FE_PHN3129_n750), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_183_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[183]), 
	.D(FE_PHN3117_n749), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_191_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[191]), 
	.D(FE_PHN3145_n748), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_199_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[199]), 
	.D(FE_PHN1465_n747), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 plain_text_reg_207_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[207]), 
	.D(FE_PHN3150_n746), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_215_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[215]), 
	.D(FE_PHN3130_n745), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_223_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[223]), 
	.D(FE_PHN3159_n744), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_231_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[231]), 
	.D(FE_PHN3119_n743), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_239_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[239]), 
	.D(n742), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_247_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[247]), 
	.D(FE_PHN3291_n741), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_255_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[255]), 
	.D(FE_PHN1070_n740), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_6_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[6]), 
	.D(FE_PHN2854_n739), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 plain_text_reg_14_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[14]), 
	.D(n738), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_22_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[22]), 
	.D(n737), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_text_reg_30_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[30]), 
	.D(FE_PHN3347_n736), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_text_reg_38_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[38]), 
	.D(FE_PHN1911_n735), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_text_reg_46_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[46]), 
	.D(FE_PHN1898_n734), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_text_reg_54_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[54]), 
	.D(n733), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 plain_text_reg_62_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[62]), 
	.D(n732), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 plain_text_reg_70_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[70]), 
	.D(n731), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 plain_text_reg_78_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[78]), 
	.D(n730), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 plain_text_reg_86_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[86]), 
	.D(n729), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_text_reg_94_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[94]), 
	.D(n728), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_text_reg_102_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[102]), 
	.D(n727), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 plain_text_reg_110_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[110]), 
	.D(FE_PHN3306_n726), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 plain_text_reg_118_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[118]), 
	.D(FE_PHN1121_n725), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 plain_text_reg_126_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[126]), 
	.D(FE_PHN3383_n724), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_134_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[134]), 
	.D(FE_PHN3155_n723), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_142_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[142]), 
	.D(FE_PHN3118_n722), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_150_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[150]), 
	.D(FE_PHN1340_n721), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_158_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[158]), 
	.D(n720), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_166_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[166]), 
	.D(FE_PHN3115_n719), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_174_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[174]), 
	.D(FE_PHN823_n718), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 plain_text_reg_182_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[182]), 
	.D(FE_PHN3172_n717), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_190_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[190]), 
	.D(FE_PHN3168_n716), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_text_reg_198_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[198]), 
	.D(FE_PHN3138_n715), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 plain_text_reg_206_ (.RN(reset_n), 
	.Q(plain_text[206]), 
	.D(FE_PHN3140_n714), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 plain_text_reg_214_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[214]), 
	.D(FE_PHN3144_n713), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 plain_text_reg_222_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[222]), 
	.D(FE_PHN3158_n712), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 plain_text_reg_230_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[230]), 
	.D(FE_PHN2851_n711), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 plain_text_reg_238_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[238]), 
	.D(FE_PHN1140_n710), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 plain_text_reg_246_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[246]), 
	.D(FE_PHN3384_n709), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_254_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[254]), 
	.D(n708), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_text_reg_5_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[5]), 
	.D(n707), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 plain_text_reg_13_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[13]), 
	.D(n706), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_21_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[21]), 
	.D(n705), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_29_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[29]), 
	.D(FE_PHN3279_n704), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_37_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[37]), 
	.D(n703), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_45_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[45]), 
	.D(n702), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_53_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[53]), 
	.D(n701), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_text_reg_61_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[61]), 
	.D(n700), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 plain_text_reg_69_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[69]), 
	.D(n699), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 plain_text_reg_77_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[77]), 
	.D(n698), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_text_reg_85_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[85]), 
	.D(n697), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_text_reg_93_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[93]), 
	.D(n696), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_text_reg_101_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[101]), 
	.D(n695), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_text_reg_109_ (.RN(FE_OFN38_reset_n), 
	.Q(plain_text[109]), 
	.D(n694), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_text_reg_117_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[117]), 
	.D(FE_PHN3361_n693), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_text_reg_125_ (.RN(FE_OFN50_reset_n), 
	.Q(plain_text[125]), 
	.D(FE_PHN1895_n692), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_text_reg_133_ (.RN(FE_OFN56_reset_n), 
	.Q(plain_text[133]), 
	.D(FE_PHN1944_n691), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_text_reg_141_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[141]), 
	.D(n690), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_text_reg_149_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[149]), 
	.D(n689), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 plain_text_reg_157_ (.RN(reset_n), 
	.Q(plain_text[157]), 
	.D(FE_PHN2881_n688), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 plain_text_reg_165_ (.RN(reset_n), 
	.Q(plain_text[165]), 
	.D(FE_PHN1939_n687), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 plain_text_reg_173_ (.RN(FE_OFN47_reset_n), 
	.Q(plain_text[173]), 
	.D(FE_PHN3381_n686), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_181_ (.RN(FE_OFN47_reset_n), 
	.Q(plain_text[181]), 
	.D(n685), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_189_ (.RN(FE_OFN47_reset_n), 
	.Q(plain_text[189]), 
	.D(n684), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_197_ (.RN(FE_OFN47_reset_n), 
	.Q(plain_text[197]), 
	.D(n683), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_205_ (.RN(FE_OFN47_reset_n), 
	.Q(plain_text[205]), 
	.D(n682), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_213_ (.RN(FE_OFN47_reset_n), 
	.Q(plain_text[213]), 
	.D(n681), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_221_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[221]), 
	.D(FE_PHN2872_n680), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_229_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[229]), 
	.D(FE_PHN1865_n679), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_237_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[237]), 
	.D(FE_PHN1927_n678), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 plain_text_reg_245_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[245]), 
	.D(FE_PHN1741_n677), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_253_ (.RN(FE_OFN58_reset_n), 
	.Q(plain_text[253]), 
	.D(FE_PHN1704_n676), 
	.CK(clk_48Mhz__L6_N20));
   DFFRHQX1 plain_text_reg_4_ (.RN(FE_OFN44_reset_n), 
	.Q(plain_text[4]), 
	.D(n675), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_text_reg_12_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[12]), 
	.D(FE_PHN2853_n674), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_text_reg_20_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[20]), 
	.D(n673), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_28_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[28]), 
	.D(n672), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_text_reg_36_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[36]), 
	.D(n671), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_44_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[44]), 
	.D(n670), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_52_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[52]), 
	.D(FE_PHN2866_n669), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_60_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[60]), 
	.D(FE_PHN1072_n668), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_68_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[68]), 
	.D(n667), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_76_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[76]), 
	.D(n666), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_84_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[84]), 
	.D(n665), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_92_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[92]), 
	.D(n664), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_100_ (.RN(FE_OFN51_reset_n), 
	.Q(plain_text[100]), 
	.D(n663), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_108_ (.RN(FE_OFN38_reset_n), 
	.Q(plain_text[108]), 
	.D(n662), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_116_ (.RN(FE_OFN38_reset_n), 
	.Q(plain_text[116]), 
	.D(FE_PHN3257_n661), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_124_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[124]), 
	.D(FE_PHN1934_n660), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_132_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[132]), 
	.D(FE_PHN1212_n659), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 plain_text_reg_140_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[140]), 
	.D(FE_PHN3370_n658), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_text_reg_148_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[148]), 
	.D(n657), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_text_reg_156_ (.RN(reset_n), 
	.Q(plain_text[156]), 
	.D(n656), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_text_reg_164_ (.RN(reset_n), 
	.Q(plain_text[164]), 
	.D(n655), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_text_reg_172_ (.RN(reset_n), 
	.Q(plain_text[172]), 
	.D(n654), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_text_reg_180_ (.RN(FE_OFN47_reset_n), 
	.Q(plain_text[180]), 
	.D(FE_PHN1914_n653), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_188_ (.RN(FE_OFN47_reset_n), 
	.Q(plain_text[188]), 
	.D(n652), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_196_ (.RN(FE_OFN47_reset_n), 
	.Q(plain_text[196]), 
	.D(FE_PHN2859_n651), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 plain_text_reg_204_ (.RN(FE_OFN47_reset_n), 
	.Q(plain_text[204]), 
	.D(n650), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_212_ (.RN(FE_OFN47_reset_n), 
	.Q(plain_text[212]), 
	.D(FE_PHN1918_n649), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_220_ (.RN(FE_OFN47_reset_n), 
	.Q(plain_text[220]), 
	.D(n648), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_228_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[228]), 
	.D(n647), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_236_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[236]), 
	.D(n646), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_244_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[244]), 
	.D(FE_PHN3264_n645), 
	.CK(clk_48Mhz__L6_N20));
   DFFRHQX1 plain_text_reg_252_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[252]), 
	.D(FE_PHN1061_n644), 
	.CK(clk_48Mhz__L6_N20));
   DFFRHQX1 plain_text_reg_3_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[3]), 
	.D(n643), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 plain_text_reg_11_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_text[11]), 
	.D(n642), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_text_reg_19_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[19]), 
	.D(FE_PHN3142_n641), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_text_reg_27_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[27]), 
	.D(FE_PHN3111_n640), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_text_reg_35_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[35]), 
	.D(FE_PHN1090_n639), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_text_reg_43_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[43]), 
	.D(FE_PHN3380_n638), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_51_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[51]), 
	.D(n637), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_59_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[59]), 
	.D(FE_PHN2858_n636), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_text_reg_67_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[67]), 
	.D(FE_PHN1929_n635), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_75_ (.RN(FE_OFN49_reset_n), 
	.Q(plain_text[75]), 
	.D(FE_PHN1926_n634), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_83_ (.RN(FE_OFN49_reset_n), 
	.Q(plain_text[83]), 
	.D(n633), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_91_ (.RN(FE_OFN49_reset_n), 
	.Q(plain_text[91]), 
	.D(n632), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_99_ (.RN(FE_OFN38_reset_n), 
	.Q(plain_text[99]), 
	.D(n631), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_107_ (.RN(FE_OFN49_reset_n), 
	.Q(plain_text[107]), 
	.D(n630), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_115_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[115]), 
	.D(n629), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_123_ (.RN(FE_OFN52_reset_n), 
	.Q(plain_text[123]), 
	.D(n628), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_text_reg_131_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[131]), 
	.D(n627), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 plain_text_reg_139_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[139]), 
	.D(FE_PHN2883_n626), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 plain_text_reg_147_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[147]), 
	.D(FE_PHN1198_n625), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 plain_text_reg_155_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[155]), 
	.D(FE_PHN3387_n624), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_text_reg_163_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[163]), 
	.D(n623), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_text_reg_171_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[171]), 
	.D(n622), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_text_reg_179_ (.RN(FE_OFN58_reset_n), 
	.Q(plain_text[179]), 
	.D(n621), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_text_reg_187_ (.RN(FE_OFN58_reset_n), 
	.Q(plain_text[187]), 
	.D(FE_PHN3385_n620), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 plain_text_reg_195_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[195]), 
	.D(FE_PHN1936_n619), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_203_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[203]), 
	.D(FE_PHN1923_n618), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_211_ (.RN(FE_OFN58_reset_n), 
	.Q(plain_text[211]), 
	.D(FE_PHN3352_n617), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_219_ (.RN(FE_OFN58_reset_n), 
	.Q(plain_text[219]), 
	.D(FE_PHN1842_n616), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_227_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[227]), 
	.D(FE_PHN1949_n615), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_235_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[235]), 
	.D(n614), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_text_reg_243_ (.RN(FE_OFN58_reset_n), 
	.Q(plain_text[243]), 
	.D(FE_PHN1928_n613), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 plain_text_reg_251_ (.RN(FE_OFN58_reset_n), 
	.Q(plain_text[251]), 
	.D(FE_PHN3300_n612), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 plain_text_reg_2_ (.RN(reset_n), 
	.Q(plain_text[2]), 
	.D(n611), 
	.CK(clk_48Mhz__L6_N25));
   DFFRHQX1 plain_text_reg_10_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[10]), 
	.D(n610), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 plain_text_reg_18_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[18]), 
	.D(FE_PHN1186_n609), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 plain_text_reg_26_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[26]), 
	.D(FE_PHN3368_n608), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_text_reg_34_ (.RN(FE_OFN56_reset_n), 
	.Q(plain_text[34]), 
	.D(n607), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_text_reg_42_ (.RN(FE_OFN56_reset_n), 
	.Q(plain_text[42]), 
	.D(FE_PHN3199_n606), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_text_reg_50_ (.RN(FE_OFN39_reset_n), 
	.Q(plain_text[50]), 
	.D(FE_PHN3366_n605), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_text_reg_58_ (.RN(FE_OFN56_reset_n), 
	.Q(plain_text[58]), 
	.D(n604), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_text_reg_66_ (.RN(FE_OFN56_reset_n), 
	.Q(plain_text[66]), 
	.D(n603), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_text_reg_74_ (.RN(FE_OFN56_reset_n), 
	.Q(plain_text[74]), 
	.D(n602), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_text_reg_82_ (.RN(FE_OFN56_reset_n), 
	.Q(plain_text[82]), 
	.D(n601), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_text_reg_90_ (.RN(FE_OFN39_reset_n), 
	.Q(plain_text[90]), 
	.D(n600), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_text_reg_98_ (.RN(FE_OFN39_reset_n), 
	.Q(plain_text[98]), 
	.D(n599), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_text_reg_106_ (.RN(FE_OFN39_reset_n), 
	.Q(plain_text[106]), 
	.D(n598), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_text_reg_114_ (.RN(FE_OFN39_reset_n), 
	.Q(plain_text[114]), 
	.D(n597), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 plain_text_reg_122_ (.RN(FE_OFN55_reset_n), 
	.Q(plain_text[122]), 
	.D(n596), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_text_reg_130_ (.RN(FE_OFN39_reset_n), 
	.Q(plain_text[130]), 
	.D(n595), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_text_reg_138_ (.RN(FE_OFN39_reset_n), 
	.Q(plain_text[138]), 
	.D(n594), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_text_reg_146_ (.RN(FE_OFN39_reset_n), 
	.Q(plain_text[146]), 
	.D(FE_PHN2886_n593), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_text_reg_154_ (.RN(FE_OFN56_reset_n), 
	.Q(plain_text[154]), 
	.D(FE_PHN1909_n592), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_text_reg_162_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[162]), 
	.D(FE_PHN1947_n591), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_text_reg_170_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[170]), 
	.D(n590), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_text_reg_178_ (.RN(FE_OFN58_reset_n), 
	.Q(plain_text[178]), 
	.D(n589), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_text_reg_186_ (.RN(FE_OFN58_reset_n), 
	.Q(plain_text[186]), 
	.D(n588), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_194_ (.RN(FE_OFN58_reset_n), 
	.Q(plain_text[194]), 
	.D(n587), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_202_ (.RN(FE_OFN58_reset_n), 
	.Q(plain_text[202]), 
	.D(n586), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_210_ (.RN(FE_OFN58_reset_n), 
	.Q(plain_text[210]), 
	.D(n585), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_text_reg_218_ (.RN(FE_OFN58_reset_n), 
	.Q(plain_text[218]), 
	.D(FE_PHN3374_n584), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 plain_text_reg_226_ (.RN(FE_OFN58_reset_n), 
	.Q(plain_text[226]), 
	.D(FE_PHN1920_n583), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 plain_text_reg_234_ (.RN(FE_OFN58_reset_n), 
	.Q(plain_text[234]), 
	.D(FE_PHN3364_n582), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_text_reg_242_ (.RN(FE_OFN58_reset_n), 
	.Q(plain_text[242]), 
	.D(FE_PHN1875_n581), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_text_reg_250_ (.RN(FE_OFN58_reset_n), 
	.Q(plain_text[250]), 
	.D(FE_PHN1815_n580), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 plain_text_reg_1_ (.RN(reset_n), 
	.Q(plain_text[1]), 
	.D(n579), 
	.CK(clk_48Mhz__L6_N28));
   DFFRHQX1 plain_text_reg_9_ (.RN(FE_OFN44_reset_n), 
	.Q(plain_text[9]), 
	.D(n578), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_text_reg_17_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[17]), 
	.D(n577), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_text_reg_25_ (.RN(FE_OFN49_reset_n), 
	.Q(plain_text[25]), 
	.D(n576), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_text_reg_33_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[33]), 
	.D(FE_PHN2889_n575), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 plain_text_reg_41_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[41]), 
	.D(FE_PHN1753_n574), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_text_reg_49_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[49]), 
	.D(FE_PHN1915_n573), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 plain_text_reg_57_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[57]), 
	.D(n572), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_text_reg_65_ (.RN(FE_OFN43_reset_n), 
	.Q(plain_text[65]), 
	.D(n571), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_text_reg_73_ (.RN(FE_OFN49_reset_n), 
	.Q(plain_text[73]), 
	.D(n570), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_text_reg_81_ (.RN(FE_OFN49_reset_n), 
	.Q(plain_text[81]), 
	.D(n569), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_text_reg_89_ (.RN(FE_OFN49_reset_n), 
	.Q(plain_text[89]), 
	.D(n568), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_text_reg_97_ (.RN(FE_OFN49_reset_n), 
	.Q(plain_text[97]), 
	.D(n567), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_text_reg_105_ (.RN(FE_OFN44_reset_n), 
	.Q(plain_text[105]), 
	.D(n566), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_text_reg_113_ (.RN(FE_OFN44_reset_n), 
	.Q(plain_text[113]), 
	.D(n565), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_text_reg_121_ (.RN(FE_OFN44_reset_n), 
	.Q(plain_text[121]), 
	.D(n564), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_text_reg_129_ (.RN(FE_OFN44_reset_n), 
	.Q(plain_text[129]), 
	.D(n563), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 plain_text_reg_137_ (.RN(FE_OFN44_reset_n), 
	.Q(plain_text[137]), 
	.D(FE_PHN3113_n562), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 plain_text_reg_145_ (.RN(FE_OFN44_reset_n), 
	.Q(plain_text[145]), 
	.D(FE_PHN2852_n561), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 plain_text_reg_153_ (.RN(FE_OFN44_reset_n), 
	.Q(plain_text[153]), 
	.D(FE_PHN1924_n560), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_text_reg_161_ (.RN(reset_n), 
	.Q(plain_text[161]), 
	.D(FE_PHN1922_n559), 
	.CK(clk_48Mhz));
   DFFRHQX1 plain_text_reg_169_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[169]), 
	.D(FE_PHN3297_n558), 
	.CK(clk_48Mhz));
   DFFRHQX1 plain_text_reg_177_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[177]), 
	.D(FE_PHN3346_n557), 
	.CK(clk_48Mhz));
   DFFRHQX1 plain_text_reg_185_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[185]), 
	.D(FE_PHN1919_n556), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_text_reg_193_ (.RN(reset_n), 
	.Q(plain_text[193]), 
	.D(FE_PHN1931_n555), 
	.CK(clk_48Mhz));
   DFFRHQX1 plain_text_reg_201_ (.RN(reset_n), 
	.Q(plain_text[201]), 
	.D(FE_PHN2873_n554), 
	.CK(clk_48Mhz));
   DFFRHQX1 plain_text_reg_209_ (.RN(FE_OFN44_reset_n), 
	.Q(plain_text[209]), 
	.D(FE_PHN1845_n553), 
	.CK(clk_48Mhz));
   DFFRHQX1 plain_text_reg_217_ (.RN(reset_n), 
	.Q(plain_text[217]), 
	.D(FE_PHN1902_n552), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_text_reg_225_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[225]), 
	.D(FE_PHN2869_n551), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_text_reg_233_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[233]), 
	.D(FE_PHN1836_n550), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_text_reg_241_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[241]), 
	.D(FE_PHN1890_n549), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_text_reg_249_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[249]), 
	.D(n548), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 plain_text_reg_0_ (.RN(FE_OFN47_reset_n), 
	.Q(plain_text[0]), 
	.D(n547), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 plain_text_reg_8_ (.RN(FE_OFN40_reset_n), 
	.Q(plain_text[8]), 
	.D(FE_PHN1203_n546), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_text_reg_16_ (.RN(FE_OFN40_reset_n), 
	.Q(plain_text[16]), 
	.D(FE_PHN3375_n545), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_text_reg_24_ (.RN(FE_OFN40_reset_n), 
	.Q(plain_text[24]), 
	.D(n544), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_text_reg_32_ (.RN(FE_OFN49_reset_n), 
	.Q(plain_text[32]), 
	.D(FE_PHN3372_n543), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_text_reg_40_ (.RN(FE_OFN49_reset_n), 
	.Q(plain_text[40]), 
	.D(FE_PHN3377_n542), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_text_reg_48_ (.RN(FE_OFN49_reset_n), 
	.Q(plain_text[48]), 
	.D(n541), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_text_reg_56_ (.RN(FE_OFN40_reset_n), 
	.Q(plain_text[56]), 
	.D(n540), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_text_reg_64_ (.RN(FE_OFN44_reset_n), 
	.Q(plain_text[64]), 
	.D(FE_PHN3132_n539), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_text_reg_72_ (.RN(FE_OFN40_reset_n), 
	.Q(plain_text[72]), 
	.D(FE_PHN3109_n538), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_text_reg_80_ (.RN(FE_OFN40_reset_n), 
	.Q(plain_text[80]), 
	.D(FE_PHN3123_n537), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_text_reg_88_ (.RN(FE_OFN40_reset_n), 
	.Q(plain_text[88]), 
	.D(n536), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_text_reg_96_ (.RN(FE_OFN40_reset_n), 
	.Q(plain_text[96]), 
	.D(n535), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_text_reg_104_ (.RN(FE_OFN44_reset_n), 
	.Q(plain_text[104]), 
	.D(n534), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_text_reg_112_ (.RN(FE_OFN44_reset_n), 
	.Q(plain_text[112]), 
	.D(n533), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_text_reg_120_ (.RN(FE_OFN44_reset_n), 
	.Q(plain_text[120]), 
	.D(n532), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_text_reg_128_ (.RN(FE_OFN44_reset_n), 
	.Q(plain_text[128]), 
	.D(n531), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 plain_text_reg_136_ (.RN(FE_OFN44_reset_n), 
	.Q(plain_text[136]), 
	.D(FE_PHN3122_n530), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_text_reg_144_ (.RN(FE_OFN44_reset_n), 
	.Q(plain_text[144]), 
	.D(FE_PHN1900_n529), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_text_reg_152_ (.RN(FE_OFN44_reset_n), 
	.Q(plain_text[152]), 
	.D(FE_PHN1938_n528), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_text_reg_160_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[160]), 
	.D(FE_PHN1912_n527), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_text_reg_168_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[168]), 
	.D(FE_PHN1932_n526), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_text_reg_176_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[176]), 
	.D(FE_PHN3134_n525), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_text_reg_184_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[184]), 
	.D(FE_PHN1886_n524), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_text_reg_192_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[192]), 
	.D(FE_PHN1933_n523), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_text_reg_200_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[200]), 
	.D(FE_PHN3286_n522), 
	.CK(clk_48Mhz));
   DFFRHQX1 plain_text_reg_208_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[208]), 
	.D(n521), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_text_reg_216_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[216]), 
	.D(n520), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_text_reg_224_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[224]), 
	.D(FE_PHN3357_n519), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_text_reg_232_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[232]), 
	.D(FE_PHN1903_n518), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_text_reg_240_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[240]), 
	.D(FE_PHN1946_n517), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_text_reg_248_ (.RN(FE_OFN45_reset_n), 
	.Q(plain_text[248]), 
	.D(FE_PHN5232_n516), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_247_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN659_Din_247_), 
	.D(FE_PHN2986_n507), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_key_out_reg_246_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN522_Din_246_), 
	.D(FE_PHN3580_n506), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_key_out_reg_245_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN476_Din_245_), 
	.D(FE_PHN3026_n505), 
	.CK(clk_48Mhz__L6_N20));
   DFFRHQX1 plain_key_out_reg_244_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN649_Din_244_), 
	.D(FE_PHN3055_n504), 
	.CK(clk_48Mhz__L6_N20));
   DFFRHQX1 plain_key_out_reg_243_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN486_Din_243_), 
	.D(FE_PHN3517_n503), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 plain_key_out_reg_242_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN474_Din_242_), 
	.D(FE_PHN5158_n502), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 plain_key_out_reg_241_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN648_Din_241_), 
	.D(FE_PHN3018_n501), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_key_out_reg_240_ (.RN(FE_OFN44_reset_n), 
	.Q(FE_PHN453_Din_240_), 
	.D(FE_PHN3445_n500), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_key_out_reg_239_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN480_Din_239_), 
	.D(FE_PHN3470_n499), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_key_out_reg_238_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN459_Din_238_), 
	.D(FE_PHN1825_n498), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_key_out_reg_237_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN652_Din_237_), 
	.D(FE_PHN3049_n497), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 plain_key_out_reg_236_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN517_Din_236_), 
	.D(FE_PHN3504_n496), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_key_out_reg_235_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN477_Din_235_), 
	.D(FE_PHN2997_n495), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_key_out_reg_234_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN490_Din_234_), 
	.D(FE_PHN3014_n494), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_key_out_reg_233_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN498_Din_233_), 
	.D(FE_PHN3047_n493), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_key_out_reg_232_ (.RN(FE_OFN44_reset_n), 
	.Q(FE_PHN456_Din_232_), 
	.D(FE_PHN2996_n492), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_key_out_reg_231_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN516_Din_231_), 
	.D(FE_PHN3405_n491), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_key_out_reg_230_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN483_Din_230_), 
	.D(FE_PHN3394_n490), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 plain_key_out_reg_229_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN499_Din_229_), 
	.D(FE_PHN3036_n489), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_key_out_reg_228_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN524_Din_228_), 
	.D(FE_PHN3582_n488), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_key_out_reg_227_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN653_Din_227_), 
	.D(FE_PHN3056_n487), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 plain_key_out_reg_226_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN520_Din_226_), 
	.D(FE_PHN1407_n486), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 plain_key_out_reg_225_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN663_Din_225_), 
	.D(FE_PHN3518_n485), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_key_out_reg_224_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN492_Din_224_), 
	.D(FE_PHN3046_n484), 
	.CK(clk_48Mhz));
   DFFRHQX1 plain_key_out_reg_223_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN475_Din_223_), 
	.D(FE_PHN3443_n483), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_key_out_reg_222_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN501_Din_222_), 
	.D(FE_PHN3498_n482), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_key_out_reg_221_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN651_Din_221_), 
	.D(FE_PHN3070_n481), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_key_out_reg_220_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN654_Din_220_), 
	.D(FE_PHN3497_n480), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_key_out_reg_219_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN532_Din_219_), 
	.D(FE_PHN3078_n479), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_key_out_reg_218_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN514_Din_218_), 
	.D(FE_PHN3071_n478), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 plain_key_out_reg_217_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN500_Din_217_), 
	.D(FE_PHN3514_n477), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_key_out_reg_216_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN464_Din_216_), 
	.D(FE_PHN3462_n476), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_key_out_reg_215_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_key_out[215]), 
	.D(FE_PHN1431_n475), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_key_out_reg_214_ (.RN(FE_OFN42_reset_n), 
	.Q(plain_key_out[214]), 
	.D(FE_PHN2794_n474), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_key_out_reg_213_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN507_Din_213_), 
	.D(FE_PHN3494_n473), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_key_out_reg_212_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN657_Din_212_), 
	.D(FE_PHN3574_n472), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_key_out_reg_211_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN670_Din_211_), 
	.D(FE_PHN3035_n471), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_key_out_reg_210_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN526_Din_210_), 
	.D(FE_PHN3598_n470), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 plain_key_out_reg_209_ (.RN(FE_OFN44_reset_n), 
	.Q(FE_PHN455_Din_209_), 
	.D(FE_PHN2962_n469), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_key_out_reg_208_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN662_Din_208_), 
	.D(FE_PHN3554_n468), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_key_out_reg_207_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN469_Din_207_), 
	.D(FE_PHN3397_n467), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_key_out_reg_206_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN470_Din_206_), 
	.D(FE_PHN3395_n466), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 plain_key_out_reg_205_ (.RN(FE_OFN47_reset_n), 
	.Q(FE_PHN497_Din_205_), 
	.D(FE_PHN3478_n465), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_key_out_reg_204_ (.RN(FE_OFN47_reset_n), 
	.Q(FE_PHN509_Din_204_), 
	.D(FE_PHN3060_n464), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_key_out_reg_203_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN513_Din_203_), 
	.D(FE_PHN3534_n463), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_key_out_reg_202_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN525_Din_202_), 
	.D(FE_PHN3561_n462), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_key_out_reg_201_ (.RN(FE_OFN44_reset_n), 
	.Q(FE_PHN467_Din_201_), 
	.D(FE_PHN3439_n461), 
	.CK(clk_48Mhz));
   DFFRHQX1 plain_key_out_reg_200_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN512_Din_200_), 
	.D(FE_PHN3545_n460), 
	.CK(clk_48Mhz));
   DFFRHQX1 plain_key_out_reg_199_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN489_Din_199_), 
	.D(FE_PHN1154_n459), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 plain_key_out_reg_198_ (.RN(reset_n), 
	.Q(FE_PHN454_Din_198_), 
	.D(FE_PHN3392_n458), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 plain_key_out_reg_197_ (.RN(FE_OFN47_reset_n), 
	.Q(FE_PHN639_Din_197_), 
	.D(FE_PHN2928_n457), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 plain_key_out_reg_196_ (.RN(FE_OFN47_reset_n), 
	.Q(FE_PHN494_Din_196_), 
	.D(FE_PHN1356_n456), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 plain_key_out_reg_195_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN508_Din_195_), 
	.D(FE_PHN3059_n455), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 plain_key_out_reg_194_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN487_Din_194_), 
	.D(FE_PHN3499_n454), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_key_out_reg_193_ (.RN(reset_n), 
	.Q(FE_PHN479_Din_193_), 
	.D(FE_PHN3455_n453), 
	.CK(clk_48Mhz));
   DFFRHQX1 plain_key_out_reg_192_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN478_Din_192_), 
	.D(FE_PHN3493_n452), 
	.CK(clk_48Mhz));
   DFFRHQX1 plain_key_out_reg_191_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN641_Din_191_), 
	.D(FE_PHN2931_n451), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 plain_key_out_reg_190_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN481_Din_190_), 
	.D(FE_PHN3495_n450), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_key_out_reg_189_ (.RN(FE_OFN47_reset_n), 
	.Q(FE_PHN529_Din_189_), 
	.D(FE_PHN3568_n449), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_key_out_reg_188_ (.RN(FE_OFN47_reset_n), 
	.Q(FE_PHN665_Din_188_), 
	.D(FE_PHN3571_n448), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_key_out_reg_187_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN527_Din_187_), 
	.D(FE_PHN3076_n447), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 plain_key_out_reg_186_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN668_Din_186_), 
	.D(FE_PHN3544_n446), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 plain_key_out_reg_185_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN519_Din_185_), 
	.D(FE_PHN3069_n445), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_key_out_reg_184_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN502_Din_184_), 
	.D(FE_PHN3053_n444), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 plain_key_out_reg_183_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN680_Din_183_), 
	.D(FE_PHN1437_n443), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_key_out_reg_182_ (.RN(FE_OFN44_reset_n), 
	.Q(FE_PHN679_Din_182_), 
	.D(FE_PHN3603_n442), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_key_out_reg_181_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN661_Din_181_), 
	.D(FE_PHN3508_n441), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_key_out_reg_180_ (.RN(FE_OFN47_reset_n), 
	.Q(FE_PHN666_Din_180_), 
	.D(FE_PHN3492_n440), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_key_out_reg_179_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN504_Din_179_), 
	.D(FE_PHN3558_n439), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 plain_key_out_reg_178_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN506_Din_178_), 
	.D(FE_PHN3539_n438), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 plain_key_out_reg_177_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN510_Din_177_), 
	.D(FE_PHN3072_n437), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_key_out_reg_176_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN485_Din_176_), 
	.D(FE_PHN3058_n436), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_key_out_reg_175_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN447_Din_175_), 
	.D(FE_PHN3393_n435), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_key_out_reg_174_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN472_Din_174_), 
	.D(FE_PHN1128_n434), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 plain_key_out_reg_173_ (.RN(FE_OFN47_reset_n), 
	.Q(FE_PHN496_Din_173_), 
	.D(FE_PHN3511_n433), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_key_out_reg_172_ (.RN(FE_OFN47_reset_n), 
	.Q(FE_PHN452_Din_172_), 
	.D(FE_PHN2967_n432), 
	.CK(clk_48Mhz__L6_N27));
   DFFRHQX1 plain_key_out_reg_171_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN468_Din_171_), 
	.D(FE_PHN3441_n431), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_key_out_reg_170_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN463_Din_170_), 
	.D(FE_PHN3440_n430), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_key_out_reg_169_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN484_Din_169_), 
	.D(FE_PHN3468_n429), 
	.CK(clk_48Mhz));
   DFFRHQX1 plain_key_out_reg_168_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN488_Din_168_), 
	.D(FE_PHN3471_n428), 
	.CK(clk_48Mhz));
   DFFRHQX1 plain_key_out_reg_167_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN637_Din_167_), 
	.D(FE_PHN711_n427), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 plain_key_out_reg_166_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN644_Din_166_), 
	.D(FE_PHN2815_n426), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 plain_key_out_reg_165_ (.RN(reset_n), 
	.Q(FE_PHN465_Din_165_), 
	.D(FE_PHN1330_n425), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 plain_key_out_reg_164_ (.RN(reset_n), 
	.Q(FE_PHN643_Din_164_), 
	.D(FE_PHN2975_n424), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 plain_key_out_reg_163_ (.RN(reset_n), 
	.Q(FE_PHN493_Din_163_), 
	.D(FE_PHN1357_n423), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 plain_key_out_reg_162_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN495_Din_162_), 
	.D(FE_PHN3028_n422), 
	.CK(clk_48Mhz__L6_N29));
   DFFRHQX1 plain_key_out_reg_161_ (.RN(reset_n), 
	.Q(FE_PHN450_Din_161_), 
	.D(FE_PHN3460_n421), 
	.CK(clk_48Mhz));
   DFFRHQX1 plain_key_out_reg_160_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN523_Din_160_), 
	.D(FE_PHN3073_n420), 
	.CK(clk_48Mhz));
   DFFRHQX1 plain_key_out_reg_159_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN667_Din_159_), 
	.D(FE_PHN3401_n419), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_key_out_reg_158_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN677_Din_158_), 
	.D(FE_PHN3399_n418), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_key_out_reg_157_ (.RN(FE_OFN47_reset_n), 
	.Q(FE_PHN676_Din_157_), 
	.D(FE_PHN3602_n417), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_key_out_reg_156_ (.RN(FE_OFN47_reset_n), 
	.Q(FE_PHN672_Din_156_), 
	.D(FE_PHN3549_n416), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_key_out_reg_155_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN675_Din_155_), 
	.D(FE_PHN3570_n415), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_key_out_reg_154_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN530_Din_154_), 
	.D(FE_PHN3077_n414), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_key_out_reg_153_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN518_Din_153_), 
	.D(FE_PHN3068_n413), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_key_out_reg_152_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN491_Din_152_), 
	.D(FE_PHN3062_n412), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_key_out_reg_151_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN660_Din_151_), 
	.D(FE_PHN3396_n411), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_key_out_reg_150_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN656_Din_150_), 
	.D(FE_PHN3402_n410), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_key_out_reg_149_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN671_Din_149_), 
	.D(FE_PHN3590_n409), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_key_out_reg_148_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN673_Din_148_), 
	.D(FE_PHN2963_n408), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 plain_key_out_reg_147_ (.RN(FE_OFN39_reset_n), 
	.Q(FE_PHN674_Din_147_), 
	.D(FE_PHN3600_n407), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_key_out_reg_146_ (.RN(FE_OFN39_reset_n), 
	.Q(FE_PHN669_Din_146_), 
	.D(FE_PHN3555_n406), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_key_out_reg_145_ (.RN(FE_OFN44_reset_n), 
	.Q(FE_PHN471_Din_145_), 
	.D(FE_PHN3513_n405), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_key_out_reg_144_ (.RN(FE_OFN44_reset_n), 
	.Q(FE_PHN466_Din_144_), 
	.D(FE_PHN2974_n404), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_key_out_reg_143_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN460_Din_143_), 
	.D(FE_PHN3447_n403), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_key_out_reg_142_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN503_Din_142_), 
	.D(FE_PHN3022_n402), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_key_out_reg_141_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN511_Din_141_), 
	.D(FE_PHN3550_n401), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_key_out_reg_140_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN655_Din_140_), 
	.D(FE_PHN3506_n400), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_key_out_reg_139_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN531_Din_139_), 
	.D(FE_PHN3604_n399), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_key_out_reg_138_ (.RN(FE_OFN39_reset_n), 
	.Q(FE_PHN473_Din_138_), 
	.D(FE_PHN3442_n398), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_key_out_reg_137_ (.RN(FE_OFN44_reset_n), 
	.Q(FE_PHN448_Din_137_), 
	.D(FE_PHN3436_n397), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 plain_key_out_reg_136_ (.RN(FE_OFN44_reset_n), 
	.Q(FE_PHN461_Din_136_), 
	.D(FE_PHN3021_n396), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 plain_key_out_reg_135_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN482_Din_135_), 
	.D(FE_PHN1136_n395), 
	.CK(clk_48Mhz__L6_N2));
   DFFRHQX1 plain_key_out_reg_134_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN515_Din_134_), 
	.D(FE_PHN3529_n394), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_key_out_reg_133_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN451_Din_133_), 
	.D(FE_PHN3466_n393), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_key_out_reg_132_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN449_Din_132_), 
	.D(FE_PHN3454_n392), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_key_out_reg_131_ (.RN(reset_n), 
	.Q(FE_PHN458_Din_131_), 
	.D(FE_PHN3451_n391), 
	.CK(clk_48Mhz__L6_N35));
   DFFRHQX1 plain_key_out_reg_130_ (.RN(FE_OFN56_reset_n), 
	.Q(FE_PHN521_Din_130_), 
	.D(FE_PHN3537_n390), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_key_out_reg_129_ (.RN(FE_OFN44_reset_n), 
	.Q(FE_PHN457_Din_129_), 
	.D(FE_PHN3457_n389), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 plain_key_out_reg_128_ (.RN(FE_OFN44_reset_n), 
	.Q(FE_PHN462_Din_128_), 
	.D(FE_PHN3448_n388), 
	.CK(clk_48Mhz__L6_N4));
   DFFRHQX1 plain_key_out_reg_255_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN647_Din_255_), 
	.D(FE_PHN3050_n515), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_key_out_reg_254_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN640_Din_254_), 
	.D(FE_PHN2938_n514), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_key_out_reg_253_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN642_Din_253_), 
	.D(FE_PHN2934_n513), 
	.CK(clk_48Mhz__L6_N20));
   DFFRHQX1 plain_key_out_reg_252_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN658_Din_252_), 
	.D(FE_PHN2937_n512), 
	.CK(clk_48Mhz__L6_N20));
   DFFRHQX1 plain_key_out_reg_251_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN645_Din_251_), 
	.D(FE_PHN2939_n511), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 plain_key_out_reg_250_ (.RN(FE_OFN58_reset_n), 
	.Q(FE_PHN664_Din_250_), 
	.D(FE_PHN2940_n510), 
	.CK(clk_48Mhz__L6_N15));
   DFFRHQX1 plain_key_out_reg_249_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN650_Din_249_), 
	.D(FE_PHN2924_n509), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_key_out_reg_248_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN446_Din_248_), 
	.D(FE_PHN1319_n508), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_119_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN1990_Din_119_), 
	.D(FE_PHN3500_n379), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_key_out_reg_118_ (.RN(FE_OFN38_reset_n), 
	.Q(FE_PHN1995_Din_118_), 
	.D(FE_PHN3575_n378), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 plain_key_out_reg_117_ (.RN(FE_OFN38_reset_n), 
	.Q(FE_PHN1950_Din_117_), 
	.D(FE_PHN3064_n377), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_key_out_reg_116_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN1973_Din_116_), 
	.D(FE_PHN3067_n376), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_115_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN1985_Din_115_), 
	.D(FE_PHN3531_n375), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_114_ (.RN(FE_OFN39_reset_n), 
	.Q(FE_PHN1278_Din_114_), 
	.D(FE_PHN3572_n374), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 plain_key_out_reg_113_ (.RN(FE_OFN44_reset_n), 
	.Q(FE_PHN1994_Din_113_), 
	.D(FE_PHN3472_n373), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_112_ (.RN(FE_OFN40_reset_n), 
	.Q(FE_PHN1999_Din_112_), 
	.D(FE_PHN3573_n372), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_key_out_reg_111_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN1986_Din_111_), 
	.D(FE_PHN3516_n371), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_key_out_reg_110_ (.RN(FE_OFN38_reset_n), 
	.Q(FE_PHN1984_Din_110_), 
	.D(FE_PHN3039_n370), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 plain_key_out_reg_109_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN1948_Din_109_), 
	.D(FE_PHN3553_n369), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_key_out_reg_108_ (.RN(FE_OFN38_reset_n), 
	.Q(FE_PHN1955_Din_108_), 
	.D(FE_PHN3459_n368), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_107_ (.RN(FE_OFN38_reset_n), 
	.Q(FE_PHN1967_Din_107_), 
	.D(FE_PHN3579_n367), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_106_ (.RN(FE_OFN55_reset_n), 
	.Q(FE_PHN1282_Din_106_), 
	.D(FE_PHN3526_n366), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 plain_key_out_reg_105_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN1981_Din_105_), 
	.D(FE_PHN3541_n365), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_104_ (.RN(FE_OFN40_reset_n), 
	.Q(FE_PHN1910_Din_104_), 
	.D(FE_PHN3487_n364), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_key_out_reg_103_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN1925_Din_103_), 
	.D(FE_PHN3547_n363), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_key_out_reg_102_ (.RN(FE_OFN38_reset_n), 
	.Q(FE_PHN1951_Din_102_), 
	.D(FE_PHN3523_n362), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 plain_key_out_reg_101_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN1964_Din_101_), 
	.D(FE_PHN3540_n361), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_key_out_reg_100_ (.RN(FE_OFN38_reset_n), 
	.Q(FE_PHN1971_Din_100_), 
	.D(FE_PHN3446_n360), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_99_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN1916_Din_99_), 
	.D(FE_PHN3483_n359), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_98_ (.RN(FE_OFN39_reset_n), 
	.Q(FE_PHN1274_Din_98_), 
	.D(FE_PHN3449_n358), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_key_out_reg_97_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN1937_Din_97_), 
	.D(FE_PHN3510_n357), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_96_ (.RN(FE_OFN40_reset_n), 
	.Q(FE_PHN1896_Din_96_), 
	.D(FE_PHN3458_n356), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_key_out_reg_87_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN1966_Din_87_), 
	.D(FE_PHN3484_n347), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_key_out_reg_86_ (.RN(FE_OFN38_reset_n), 
	.Q(FE_PHN1963_Din_86_), 
	.D(FE_PHN3476_n346), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_key_out_reg_85_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN1975_Din_85_), 
	.D(FE_PHN3546_n345), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_key_out_reg_84_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN1956_Din_84_), 
	.D(FE_PHN3525_n344), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_83_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN1968_Din_83_), 
	.D(FE_PHN3479_n343), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_82_ (.RN(FE_OFN39_reset_n), 
	.Q(FE_PHN1908_Din_82_), 
	.D(FE_PHN3521_n342), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_key_out_reg_81_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN1281_Din_81_), 
	.D(FE_PHN3505_n341), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_80_ (.RN(FE_OFN40_reset_n), 
	.Q(FE_PHN1291_Din_80_), 
	.D(FE_PHN3465_n340), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_key_out_reg_79_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN1276_Din_79_), 
	.D(FE_PHN3548_n339), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_key_out_reg_78_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN1943_Din_78_), 
	.D(FE_PHN3473_n338), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 plain_key_out_reg_77_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN1953_Din_77_), 
	.D(FE_PHN3532_n337), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_key_out_reg_76_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN1907_Din_76_), 
	.D(FE_PHN3450_n336), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_75_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN1913_Din_75_), 
	.D(FE_PHN3461_n335), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_74_ (.RN(FE_OFN56_reset_n), 
	.Q(FE_PHN1287_Din_74_), 
	.D(FE_PHN3512_n334), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_key_out_reg_73_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN1290_Din_73_), 
	.D(FE_PHN3564_n333), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_72_ (.RN(FE_OFN40_reset_n), 
	.Q(FE_PHN1266_Din_72_), 
	.D(FE_PHN3456_n332), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_71_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN1297_Din_71_), 
	.D(FE_PHN3566_n331), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_key_out_reg_70_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN1952_Din_70_), 
	.D(FE_PHN3533_n330), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 plain_key_out_reg_69_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN1961_Din_69_), 
	.D(FE_PHN3599_n329), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_key_out_reg_68_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN1300_Din_68_), 
	.D(FE_PHN3557_n328), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_67_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN1301_Din_67_), 
	.D(FE_PHN3061_n327), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_66_ (.RN(FE_OFN56_reset_n), 
	.Q(FE_PHN1296_Din_66_), 
	.D(FE_PHN3527_n326), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_key_out_reg_65_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN1283_Din_65_), 
	.D(FE_PHN3496_n325), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_64_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN1293_Din_64_), 
	.D(FE_PHN3501_n324), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_55_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN2920_Din_55_), 
	.D(FE_PHN1906_n315), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_key_out_reg_54_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN1977_Din_54_), 
	.D(FE_PHN3583_n314), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 plain_key_out_reg_53_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN1970_Din_53_), 
	.D(FE_PHN3432_n313), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 plain_key_out_reg_52_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN1960_Din_52_), 
	.D(FE_PHN3482_n312), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_51_ (.RN(FE_OFN40_reset_n), 
	.Q(FE_PHN1978_Din_51_), 
	.D(FE_PHN3477_n311), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_50_ (.RN(FE_OFN39_reset_n), 
	.Q(FE_PHN1286_Din_50_), 
	.D(FE_PHN3485_n310), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_key_out_reg_49_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN1275_Din_49_), 
	.D(FE_PHN3467_n309), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_48_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN1292_Din_48_), 
	.D(FE_PHN3528_n308), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_47_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN1267_Din_47_), 
	.D(FE_PHN3522_n307), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_key_out_reg_46_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN1945_Din_46_), 
	.D(FE_PHN3474_n306), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_key_out_reg_45_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN1941_Din_45_), 
	.D(FE_PHN3463_n305), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_key_out_reg_44_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN1294_Din_44_), 
	.D(FE_PHN3481_n304), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_43_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN1940_Din_43_), 
	.D(FE_PHN3520_n303), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_42_ (.RN(FE_OFN56_reset_n), 
	.Q(FE_PHN1280_Din_42_), 
	.D(FE_PHN3480_n302), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_key_out_reg_41_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN1273_Din_41_), 
	.D(FE_PHN3066_n301), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_key_out_reg_40_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN1285_Din_40_), 
	.D(FE_PHN3543_n300), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_39_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN1277_Din_39_), 
	.D(FE_PHN3438_n299), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_key_out_reg_38_ (.RN(FE_OFN38_reset_n), 
	.Q(FE_PHN1306_Din_38_), 
	.D(FE_PHN3075_n298), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_key_out_reg_37_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN1942_Din_37_), 
	.D(FE_PHN3488_n297), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_key_out_reg_36_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN1303_Din_36_), 
	.D(FE_PHN3515_n296), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_35_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN1298_Din_35_), 
	.D(FE_PHN3567_n295), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_34_ (.RN(FE_OFN56_reset_n), 
	.Q(FE_PHN1271_Din_34_), 
	.D(FE_PHN3452_n294), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 plain_key_out_reg_33_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN1260_Din_33_), 
	.D(FE_PHN3475_n293), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_key_out_reg_32_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN1270_Din_32_), 
	.D(FE_PHN3536_n292), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_23_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN2921_Din_23_), 
	.D(FE_PHN1904_n283), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_key_out_reg_22_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN1279_Din_22_), 
	.D(FE_PHN3530_n282), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_key_out_reg_21_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN2922_Din_21_), 
	.D(FE_PHN1901_n281), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_key_out_reg_20_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN1982_Din_20_), 
	.D(FE_PHN3502_n280), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_19_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN1993_Din_19_), 
	.D(FE_PHN3490_n279), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_key_out_reg_18_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN1979_Din_18_), 
	.D(FE_PHN3595_n278), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_key_out_reg_17_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN1987_Din_17_), 
	.D(FE_PHN3591_n277), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_16_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN1976_Din_16_), 
	.D(FE_PHN3507_n276), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_15_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN1980_Din_15_), 
	.D(FE_PHN3535_n275), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_key_out_reg_14_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN1269_Din_14_), 
	.D(FE_PHN3562_n274), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_key_out_reg_13_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN1983_Din_13_), 
	.D(FE_PHN3552_n273), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_key_out_reg_12_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN2923_Din_12_), 
	.D(FE_PHN1423_n272), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_key_out_reg_11_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN1988_Din_11_), 
	.D(FE_PHN3593_n271), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_key_out_reg_10_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN1954_Din_10_), 
	.D(FE_PHN3596_n270), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_key_out_reg_9_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN1272_Din_9_), 
	.D(FE_PHN3469_n269), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_8_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN1268_Din_8_), 
	.D(FE_PHN3464_n268), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_7_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN1302_Din_7_), 
	.D(FE_PHN3592_n267), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_key_out_reg_6_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN1295_Din_6_), 
	.D(FE_PHN3578_n266), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_key_out_reg_5_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN1309_Din_5_), 
	.D(FE_PHN3610_n265), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_key_out_reg_4_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN1996_Din_4_), 
	.D(FE_PHN3586_n264), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_key_out_reg_3_ (.RN(FE_OFN40_reset_n), 
	.Q(FE_PHN1305_Din_3_), 
	.D(FE_PHN3584_n263), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_key_out_reg_2_ (.RN(FE_OFN45_reset_n), 
	.Q(FE_PHN1308_Din_2_), 
	.D(FE_PHN3608_n262), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_1_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN1307_Din_1_), 
	.D(FE_PHN3606_n261), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_0_ (.RN(FE_OFN40_reset_n), 
	.Q(FE_PHN1304_Din_0_), 
	.D(FE_PHN3589_n260), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_127_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN2819_Din_127_), 
	.D(FE_PHN1935_n387), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_key_out_reg_126_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN2818_Din_126_), 
	.D(FE_PHN1435_n386), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 plain_key_out_reg_125_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN749_Din_125_), 
	.D(FE_PHN2796_n385), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 plain_key_out_reg_124_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN909_Din_124_), 
	.D(FE_PHN3080_n384), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_123_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN1213_Din_123_), 
	.D(FE_PHN3609_n383), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_122_ (.RN(FE_OFN55_reset_n), 
	.Q(FE_PHN902_Din_122_), 
	.D(FE_PHN3601_n382), 
	.CK(clk_48Mhz__L6_N21));
   DFFRHQX1 plain_key_out_reg_121_ (.RN(FE_OFN44_reset_n), 
	.Q(FE_PHN1217_Din_121_), 
	.D(FE_PHN3569_n381), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_key_out_reg_120_ (.RN(FE_OFN40_reset_n), 
	.Q(FE_PHN1459_Din_120_), 
	.D(FE_PHN3560_n380), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_key_out_reg_95_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN891_Din_95_), 
	.D(FE_PHN3542_n355), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_94_ (.RN(FE_OFN38_reset_n), 
	.Q(FE_PHN906_Din_94_), 
	.D(FE_PHN3503_n354), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 plain_key_out_reg_93_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN911_Din_93_), 
	.D(FE_PHN3563_n353), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_key_out_reg_92_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN889_Din_92_), 
	.D(FE_PHN3524_n352), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_91_ (.RN(FE_OFN38_reset_n), 
	.Q(FE_PHN900_Din_91_), 
	.D(FE_PHN3581_n351), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 plain_key_out_reg_90_ (.RN(FE_OFN39_reset_n), 
	.Q(FE_PHN897_Din_90_), 
	.D(FE_PHN3486_n350), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_key_out_reg_89_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN890_Din_89_), 
	.D(FE_PHN3538_n349), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_88_ (.RN(FE_OFN40_reset_n), 
	.Q(FE_PHN904_Din_88_), 
	.D(FE_PHN3519_n348), 
	.CK(clk_48Mhz__L6_N11));
   DFFRHQX1 plain_key_out_reg_63_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN895_Din_63_), 
	.D(FE_PHN3398_n323), 
	.CK(clk_48Mhz__L6_N9));
   DFFRHQX1 plain_key_out_reg_62_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN894_Din_62_), 
	.D(FE_PHN3453_n322), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 plain_key_out_reg_61_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN892_Din_61_), 
	.D(FE_PHN3509_n321), 
	.CK(clk_48Mhz__L6_N37));
   DFFRHQX1 plain_key_out_reg_60_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN899_Din_60_), 
	.D(FE_PHN3491_n320), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_59_ (.RN(FE_OFN40_reset_n), 
	.Q(FE_PHN901_Din_59_), 
	.D(FE_PHN3587_n319), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_58_ (.RN(FE_OFN56_reset_n), 
	.Q(FE_PHN893_Din_58_), 
	.D(FE_PHN3585_n318), 
	.CK(clk_48Mhz__L6_N14));
   DFFRHQX1 plain_key_out_reg_57_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN898_Din_57_), 
	.D(FE_PHN3556_n317), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_56_ (.RN(FE_OFN40_reset_n), 
	.Q(FE_PHN903_Din_56_), 
	.D(FE_PHN3565_n316), 
	.CK(clk_48Mhz__L6_N8));
   DFFRHQX1 plain_key_out_reg_31_ (.RN(FE_OFN51_reset_n), 
	.Q(FE_PHN2817_Din_31_), 
	.D(FE_PHN1897_n291), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_key_out_reg_30_ (.RN(FE_OFN50_reset_n), 
	.Q(FE_PHN742_Din_30_), 
	.D(FE_PHN3057_n290), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 plain_key_out_reg_29_ (.RN(FE_OFN42_reset_n), 
	.Q(FE_PHN1214_Din_29_), 
	.D(FE_PHN3551_n289), 
	.CK(clk_48Mhz__L6_N5));
   DFFRHQX1 plain_key_out_reg_28_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN1215_Din_28_), 
	.D(FE_PHN3577_n288), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 plain_key_out_reg_27_ (.RN(FE_OFN52_reset_n), 
	.Q(FE_PHN1216_Din_27_), 
	.D(FE_PHN3042_n287), 
	.CK(clk_48Mhz__L6_N6));
   DFFRHQX1 plain_key_out_reg_26_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN908_Din_26_), 
	.D(FE_PHN3489_n286), 
	.CK(clk_48Mhz__L6_N23));
   DFFRHQX1 plain_key_out_reg_25_ (.RN(FE_OFN43_reset_n), 
	.Q(FE_PHN907_Din_25_), 
	.D(FE_PHN3605_n285), 
	.CK(clk_48Mhz__L6_N40));
   DFFRHQX1 plain_key_out_reg_24_ (.RN(FE_OFN49_reset_n), 
	.Q(FE_PHN910_Din_24_), 
	.D(FE_PHN3594_n284), 
	.CK(clk_48Mhz__L6_N10));
   DFFRHQX1 pbv1_reg (.RN(FE_OFN42_reset_n), 
	.Q(pbv1), 
	.D(FE_PHN5067_pbv0), 
	.CK(clk_48Mhz__L6_N1));
   DFFRHQX1 pf1_reg (.RN(FE_OFN42_reset_n), 
	.Q(pf1), 
	.D(FE_PHN5069_pf0), 
	.CK(clk_48Mhz__L6_N1));
   DFFRHQX1 pf0_reg (.RN(FE_OFN42_reset_n), 
	.Q(pf0), 
	.D(plain_finish), 
	.CK(clk_48Mhz__L6_N1));
   DFFRHQX1 pbv0_reg (.RN(FE_OFN42_reset_n), 
	.Q(pbv0), 
	.D(plain_byte_valid), 
	.CK(clk_48Mhz__L6_N1));
   INVX1 U109 (.Y(n78), 
	.A(n171));
   INVX1 U135 (.Y(n52), 
	.A(n210));
   INVX1 U185 (.Y(n153), 
	.A(n210));
   INVX1 U203 (.Y(n171), 
	.A(FE_OFN66_n258));
   CLKINVX3 U260 (.Y(n210), 
	.A(n258));
   OAI22X1 U261 (.Y(n517), 
	.B1(n1035), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1034));
   OAI22X1 U262 (.Y(n518), 
	.B1(n1034), 
	.B0(FE_OFN63_n210), 
	.A1(n153), 
	.A0(n1033));
   OAI22X1 U263 (.Y(n519), 
	.B1(n1033), 
	.B0(FE_OFN63_n210), 
	.A1(n153), 
	.A0(n1032));
   OAI22X1 U264 (.Y(n520), 
	.B1(n1032), 
	.B0(FE_OFN63_n210), 
	.A1(n153), 
	.A0(n1031));
   OAI22X1 U265 (.Y(n521), 
	.B1(n1031), 
	.B0(FE_OFN63_n210), 
	.A1(n153), 
	.A0(n1030));
   OAI22X1 U266 (.Y(n522), 
	.B1(n1030), 
	.B0(FE_OFN63_n210), 
	.A1(n153), 
	.A0(n1029));
   OAI22X1 U267 (.Y(n523), 
	.B1(n1029), 
	.B0(FE_OFN63_n210), 
	.A1(n153), 
	.A0(n1028));
   OAI22X1 U268 (.Y(n524), 
	.B1(n1028), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1027));
   OAI22X1 U269 (.Y(n525), 
	.B1(n1027), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1026));
   OAI22X1 U270 (.Y(n526), 
	.B1(n1026), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1025));
   OAI22X1 U271 (.Y(n527), 
	.B1(n1025), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1024));
   OAI22X1 U272 (.Y(n528), 
	.B1(n1024), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1023));
   OAI22X1 U273 (.Y(n529), 
	.B1(n1023), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1022));
   OAI22X1 U274 (.Y(n530), 
	.B1(n1022), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1021));
   OAI22X1 U275 (.Y(n531), 
	.B1(n1021), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1020));
   OAI22X1 U276 (.Y(n532), 
	.B1(n1020), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1019));
   OAI22X1 U277 (.Y(n533), 
	.B1(n1019), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1018));
   OAI22X1 U278 (.Y(n534), 
	.B1(n1018), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1017));
   OAI22X1 U279 (.Y(n535), 
	.B1(n1017), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1016));
   OAI22X1 U280 (.Y(n536), 
	.B1(n1016), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1015));
   OAI22X1 U281 (.Y(n537), 
	.B1(n1015), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1014));
   OAI22X1 U282 (.Y(n538), 
	.B1(n1014), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1013));
   OAI22X1 U283 (.Y(n539), 
	.B1(n1013), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1012));
   OAI22X1 U284 (.Y(n540), 
	.B1(n1012), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1011));
   OAI22X1 U285 (.Y(n541), 
	.B1(n1011), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1010));
   OAI22X1 U286 (.Y(n542), 
	.B1(n1010), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1009));
   OAI22X1 U287 (.Y(n543), 
	.B1(n1009), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1008));
   OAI22X1 U288 (.Y(n544), 
	.B1(n1008), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1007));
   OAI22X1 U289 (.Y(n545), 
	.B1(n1007), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1006));
   OAI22X1 U290 (.Y(n546), 
	.B1(n1006), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1005));
   OAI22X1 U291 (.Y(n549), 
	.B1(n1003), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1002));
   OAI22X1 U292 (.Y(n550), 
	.B1(n1002), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1001));
   OAI22X1 U293 (.Y(n551), 
	.B1(n1001), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1000));
   OAI22X1 U294 (.Y(n552), 
	.B1(n1000), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n999));
   OAI22X1 U295 (.Y(n553), 
	.B1(n999), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n998));
   OAI22X1 U296 (.Y(n554), 
	.B1(n998), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n997));
   OAI22X1 U297 (.Y(n555), 
	.B1(n997), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n996));
   OAI22X1 U298 (.Y(n556), 
	.B1(n996), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n995));
   OAI22X1 U299 (.Y(n557), 
	.B1(n995), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n994));
   OAI22X1 U300 (.Y(n558), 
	.B1(n994), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n993));
   OAI22X1 U301 (.Y(n559), 
	.B1(n993), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n992));
   OAI22X1 U302 (.Y(n560), 
	.B1(n992), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n991));
   OAI22X1 U303 (.Y(n561), 
	.B1(n991), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n990));
   OAI22X1 U304 (.Y(n562), 
	.B1(n990), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n989));
   OAI22X1 U305 (.Y(n563), 
	.B1(n989), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n988));
   OAI22X1 U306 (.Y(n564), 
	.B1(n988), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n987));
   OAI22X1 U307 (.Y(n565), 
	.B1(n987), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n986));
   OAI22X1 U308 (.Y(n566), 
	.B1(n986), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n985));
   OAI22X1 U309 (.Y(n567), 
	.B1(n985), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n984));
   OAI22X1 U310 (.Y(n568), 
	.B1(n984), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n983));
   OAI22X1 U311 (.Y(n569), 
	.B1(n983), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n982));
   OAI22X1 U312 (.Y(n570), 
	.B1(n982), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n981));
   OAI22X1 U313 (.Y(n571), 
	.B1(n981), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n980));
   OAI22X1 U314 (.Y(n572), 
	.B1(n980), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n979));
   OAI22X1 U315 (.Y(n573), 
	.B1(n979), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n978));
   OAI22X1 U316 (.Y(n574), 
	.B1(n978), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n977));
   OAI22X1 U317 (.Y(n575), 
	.B1(n977), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n976));
   OAI22X1 U318 (.Y(n576), 
	.B1(n976), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n975));
   OAI22X1 U319 (.Y(n577), 
	.B1(n975), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n974));
   OAI22X1 U320 (.Y(n578), 
	.B1(n974), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n973));
   OAI22X1 U321 (.Y(n581), 
	.B1(n971), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n970));
   OAI22X1 U322 (.Y(n582), 
	.B1(n970), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n969));
   OAI22X1 U323 (.Y(n583), 
	.B1(n969), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n968));
   OAI22X1 U324 (.Y(n584), 
	.B1(n968), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n967));
   OAI22X1 U325 (.Y(n585), 
	.B1(n967), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n966));
   OAI22X1 U326 (.Y(n586), 
	.B1(n966), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n965));
   OAI22X1 U327 (.Y(n587), 
	.B1(n965), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n964));
   OAI22X1 U328 (.Y(n588), 
	.B1(n964), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n963));
   OAI22X1 U329 (.Y(n589), 
	.B1(n963), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n962));
   OAI22X1 U330 (.Y(n590), 
	.B1(n962), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n961));
   OAI22X1 U331 (.Y(n591), 
	.B1(n961), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n960));
   OAI22X1 U332 (.Y(n592), 
	.B1(n960), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n959));
   OAI22X1 U333 (.Y(n593), 
	.B1(n959), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n958));
   OAI22X1 U334 (.Y(n594), 
	.B1(n958), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n957));
   OAI22X1 U335 (.Y(n595), 
	.B1(n957), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n956));
   OAI22X1 U336 (.Y(n596), 
	.B1(n956), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n955));
   OAI22X1 U337 (.Y(n597), 
	.B1(n955), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n954));
   OAI22X1 U338 (.Y(n598), 
	.B1(n954), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n953));
   OAI22X1 U339 (.Y(n599), 
	.B1(n953), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n952));
   OAI22X1 U340 (.Y(n600), 
	.B1(n952), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n951));
   OAI22X1 U341 (.Y(n601), 
	.B1(n951), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n950));
   OAI22X1 U342 (.Y(n602), 
	.B1(n950), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n949));
   OAI22X1 U343 (.Y(n603), 
	.B1(n949), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n948));
   OAI22X1 U344 (.Y(n604), 
	.B1(n948), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n947));
   OAI22X1 U345 (.Y(n605), 
	.B1(n947), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n946));
   OAI22X1 U346 (.Y(n606), 
	.B1(n946), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n945));
   OAI22X1 U347 (.Y(n607), 
	.B1(n945), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n944));
   OAI22X1 U348 (.Y(n608), 
	.B1(n944), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n943));
   OAI22X1 U349 (.Y(n609), 
	.B1(n943), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n942));
   OAI22X1 U350 (.Y(n610), 
	.B1(n942), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n941));
   OAI22X1 U351 (.Y(n613), 
	.B1(n939), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n938));
   OAI22X1 U352 (.Y(n614), 
	.B1(n938), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n937));
   OAI22X1 U353 (.Y(n615), 
	.B1(n937), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n936));
   OAI22X1 U354 (.Y(n616), 
	.B1(n936), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n935));
   OAI22X1 U355 (.Y(n617), 
	.B1(n935), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n934));
   OAI22X1 U356 (.Y(n618), 
	.B1(n934), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n933));
   OAI22X1 U357 (.Y(n619), 
	.B1(n933), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n932));
   OAI22X1 U358 (.Y(n620), 
	.B1(n932), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n931));
   OAI22X1 U359 (.Y(n621), 
	.B1(n931), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n930));
   OAI22X1 U360 (.Y(n622), 
	.B1(n930), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n929));
   OAI22X1 U361 (.Y(n623), 
	.B1(n929), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n928));
   OAI22X1 U362 (.Y(n624), 
	.B1(n928), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n927));
   OAI22X1 U363 (.Y(n625), 
	.B1(n927), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n926));
   OAI22X1 U364 (.Y(n626), 
	.B1(n926), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n925));
   OAI22X1 U365 (.Y(n627), 
	.B1(n925), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n924));
   OAI22X1 U366 (.Y(n628), 
	.B1(n924), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n923));
   OAI22X1 U367 (.Y(n629), 
	.B1(n923), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n922));
   OAI22X1 U368 (.Y(n630), 
	.B1(n922), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n921));
   OAI22X1 U369 (.Y(n631), 
	.B1(n921), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n920));
   OAI22X1 U370 (.Y(n632), 
	.B1(n920), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n919));
   OAI22X1 U371 (.Y(n633), 
	.B1(n919), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n918));
   OAI22X1 U372 (.Y(n634), 
	.B1(n918), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n917));
   OAI22X1 U373 (.Y(n635), 
	.B1(n917), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n916));
   OAI22X1 U374 (.Y(n636), 
	.B1(n916), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n915));
   OAI22X1 U375 (.Y(n637), 
	.B1(n915), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n914));
   OAI22X1 U376 (.Y(n638), 
	.B1(n914), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n913));
   OAI22X1 U377 (.Y(n639), 
	.B1(n913), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n912));
   OAI22X1 U378 (.Y(n640), 
	.B1(n912), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n911));
   OAI22X1 U379 (.Y(n641), 
	.B1(n911), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n910));
   OAI22X1 U380 (.Y(n642), 
	.B1(n910), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n909));
   OAI22X1 U381 (.Y(n645), 
	.B1(n907), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n906));
   OAI22X1 U382 (.Y(n646), 
	.B1(n906), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n905));
   OAI22X1 U383 (.Y(n647), 
	.B1(n905), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n904));
   OAI22X1 U384 (.Y(n648), 
	.B1(n904), 
	.B0(FE_OFN62_n210), 
	.A1(n78), 
	.A0(n903));
   OAI22X1 U385 (.Y(n649), 
	.B1(n903), 
	.B0(FE_OFN62_n210), 
	.A1(n78), 
	.A0(n902));
   OAI22X1 U386 (.Y(n650), 
	.B1(n902), 
	.B0(FE_OFN62_n210), 
	.A1(n78), 
	.A0(n901));
   OAI22X1 U387 (.Y(n651), 
	.B1(n901), 
	.B0(FE_OFN62_n210), 
	.A1(n78), 
	.A0(n900));
   OAI22X1 U388 (.Y(n652), 
	.B1(n900), 
	.B0(FE_OFN62_n210), 
	.A1(n78), 
	.A0(n899));
   OAI22X1 U389 (.Y(n653), 
	.B1(n899), 
	.B0(FE_OFN62_n210), 
	.A1(n78), 
	.A0(n898));
   OAI22X1 U390 (.Y(n654), 
	.B1(n898), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n897));
   OAI22X1 U391 (.Y(n655), 
	.B1(n897), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n896));
   OAI22X1 U392 (.Y(n656), 
	.B1(n896), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n895));
   OAI22X1 U393 (.Y(n657), 
	.B1(n895), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n894));
   OAI22X1 U394 (.Y(n658), 
	.B1(n894), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n893));
   OAI22X1 U395 (.Y(n659), 
	.B1(n893), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n892));
   OAI22X1 U396 (.Y(n660), 
	.B1(n892), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n891));
   OAI22X1 U397 (.Y(n661), 
	.B1(n891), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n890));
   OAI22X1 U398 (.Y(n662), 
	.B1(n890), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n889));
   OAI22X1 U399 (.Y(n663), 
	.B1(n889), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n888));
   OAI22X1 U400 (.Y(n664), 
	.B1(n888), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n887));
   OAI22X1 U401 (.Y(n665), 
	.B1(n887), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n886));
   OAI22X1 U402 (.Y(n666), 
	.B1(n886), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n885));
   OAI22X1 U403 (.Y(n667), 
	.B1(n885), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n884));
   OAI22X1 U404 (.Y(n668), 
	.B1(n884), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n883));
   OAI22X1 U405 (.Y(n669), 
	.B1(n883), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n882));
   OAI22X1 U406 (.Y(n670), 
	.B1(n882), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n881));
   OAI22X1 U407 (.Y(n671), 
	.B1(n881), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n880));
   OAI22X1 U408 (.Y(n672), 
	.B1(n880), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n879));
   OAI22X1 U409 (.Y(n673), 
	.B1(n879), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n878));
   OAI22X1 U410 (.Y(n674), 
	.B1(n878), 
	.B0(n210), 
	.A1(FE_OFN65_n258), 
	.A0(n877));
   OAI22X1 U411 (.Y(n677), 
	.B1(n875), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n874));
   OAI22X1 U412 (.Y(n678), 
	.B1(n874), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n873));
   OAI22X1 U413 (.Y(n679), 
	.B1(n873), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n872));
   OAI22X1 U414 (.Y(n680), 
	.B1(n872), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n871));
   OAI22X1 U415 (.Y(n681), 
	.B1(n871), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n870));
   OAI22X1 U416 (.Y(n682), 
	.B1(n870), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n869));
   OAI22X1 U417 (.Y(n683), 
	.B1(n869), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n868));
   OAI22X1 U418 (.Y(n684), 
	.B1(n868), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n867));
   OAI22X1 U419 (.Y(n685), 
	.B1(n867), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n866));
   OAI22X1 U420 (.Y(n686), 
	.B1(n866), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n865));
   OAI22X1 U421 (.Y(n687), 
	.B1(n865), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n864));
   OAI22X1 U422 (.Y(n688), 
	.B1(n864), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n863));
   OAI22X1 U423 (.Y(n689), 
	.B1(n863), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n862));
   OAI22X1 U424 (.Y(n690), 
	.B1(n862), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n861));
   OAI22X1 U425 (.Y(n691), 
	.B1(n861), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n860));
   OAI22X1 U426 (.Y(n692), 
	.B1(n860), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n859));
   OAI22X1 U427 (.Y(n693), 
	.B1(n859), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n858));
   OAI22X1 U428 (.Y(n694), 
	.B1(n858), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n857));
   OAI22X1 U429 (.Y(n695), 
	.B1(n857), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n856));
   OAI22X1 U430 (.Y(n696), 
	.B1(n856), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n855));
   OAI22X1 U431 (.Y(n697), 
	.B1(n855), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n854));
   OAI22X1 U432 (.Y(n698), 
	.B1(n854), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n853));
   OAI22X1 U433 (.Y(n699), 
	.B1(n853), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n852));
   OAI22X1 U434 (.Y(n700), 
	.B1(n852), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n851));
   OAI22X1 U435 (.Y(n701), 
	.B1(n851), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n850));
   OAI22X1 U436 (.Y(n702), 
	.B1(n850), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n849));
   OAI22X1 U437 (.Y(n703), 
	.B1(n849), 
	.B0(FE_OFN60_n210), 
	.A1(n52), 
	.A0(n848));
   OAI22X1 U438 (.Y(n704), 
	.B1(n848), 
	.B0(FE_OFN60_n210), 
	.A1(n52), 
	.A0(n847));
   OAI22X1 U439 (.Y(n705), 
	.B1(n847), 
	.B0(FE_OFN60_n210), 
	.A1(n52), 
	.A0(n846));
   OAI22X1 U440 (.Y(n706), 
	.B1(n846), 
	.B0(FE_OFN60_n210), 
	.A1(n52), 
	.A0(n845));
   OAI22X1 U441 (.Y(n709), 
	.B1(n843), 
	.B0(FE_OFN61_n210), 
	.A1(n52), 
	.A0(n842));
   OAI22X1 U442 (.Y(n710), 
	.B1(n842), 
	.B0(n210), 
	.A1(n52), 
	.A0(n841));
   OAI22X1 U443 (.Y(n711), 
	.B1(n841), 
	.B0(n210), 
	.A1(n52), 
	.A0(n840));
   OAI22X1 U444 (.Y(n712), 
	.B1(n840), 
	.B0(n210), 
	.A1(n52), 
	.A0(n839));
   OAI22X1 U445 (.Y(n713), 
	.B1(n839), 
	.B0(n210), 
	.A1(n52), 
	.A0(n838));
   OAI22X1 U446 (.Y(n714), 
	.B1(n838), 
	.B0(n210), 
	.A1(n52), 
	.A0(n837));
   OAI22X1 U447 (.Y(n715), 
	.B1(n837), 
	.B0(n210), 
	.A1(n52), 
	.A0(n836));
   OAI22X1 U448 (.Y(n716), 
	.B1(n836), 
	.B0(n210), 
	.A1(FE_OFN64_n258), 
	.A0(n835));
   OAI22X1 U449 (.Y(n717), 
	.B1(n835), 
	.B0(n210), 
	.A1(FE_OFN64_n258), 
	.A0(n834));
   OAI22X1 U450 (.Y(n718), 
	.B1(n834), 
	.B0(n210), 
	.A1(FE_PHN704_n258), 
	.A0(n833));
   OAI22X1 U451 (.Y(n719), 
	.B1(n833), 
	.B0(n210), 
	.A1(FE_PHN704_n258), 
	.A0(n832));
   OAI22X1 U452 (.Y(n720), 
	.B1(n832), 
	.B0(n210), 
	.A1(FE_PHN704_n258), 
	.A0(n831));
   OAI22X1 U453 (.Y(n721), 
	.B1(n831), 
	.B0(FE_OFN60_n210), 
	.A1(FE_PHN704_n258), 
	.A0(n830));
   OAI22X1 U454 (.Y(n722), 
	.B1(n830), 
	.B0(n210), 
	.A1(FE_PHN704_n258), 
	.A0(n829));
   OAI22X1 U455 (.Y(n723), 
	.B1(n829), 
	.B0(n210), 
	.A1(FE_PHN704_n258), 
	.A0(n828));
   OAI22X1 U456 (.Y(n724), 
	.B1(n828), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n827));
   OAI22X1 U457 (.Y(n725), 
	.B1(n827), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n826));
   OAI22X1 U458 (.Y(n726), 
	.B1(n826), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n825));
   OAI22X1 U459 (.Y(n727), 
	.B1(n825), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n824));
   OAI22X1 U460 (.Y(n728), 
	.B1(n824), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n823));
   OAI22X1 U461 (.Y(n729), 
	.B1(n823), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n822));
   OAI22X1 U462 (.Y(n730), 
	.B1(n822), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n821));
   OAI22X1 U463 (.Y(n731), 
	.B1(n821), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n820));
   OAI22X1 U464 (.Y(n732), 
	.B1(n820), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n819));
   OAI22X1 U465 (.Y(n733), 
	.B1(n819), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n818));
   OAI22X1 U466 (.Y(n734), 
	.B1(n818), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n817));
   OAI22X1 U467 (.Y(n735), 
	.B1(n817), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n816));
   OAI22X1 U468 (.Y(n736), 
	.B1(n816), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n815));
   OAI22X1 U469 (.Y(n737), 
	.B1(n815), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n814));
   OAI22X1 U470 (.Y(n738), 
	.B1(n814), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n813));
   OAI22X1 U471 (.Y(n741), 
	.B1(n811), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n810));
   OAI22X1 U472 (.Y(n742), 
	.B1(n810), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n809));
   OAI22X1 U473 (.Y(n743), 
	.B1(n809), 
	.B0(n210), 
	.A1(FE_OFN64_n258), 
	.A0(n808));
   OAI22X1 U474 (.Y(n744), 
	.B1(n808), 
	.B0(n210), 
	.A1(FE_OFN64_n258), 
	.A0(n807));
   OAI22X1 U475 (.Y(n745), 
	.B1(n807), 
	.B0(n210), 
	.A1(FE_OFN64_n258), 
	.A0(n806));
   OAI22X1 U476 (.Y(n746), 
	.B1(n806), 
	.B0(n210), 
	.A1(FE_OFN64_n258), 
	.A0(n805));
   OAI22X1 U477 (.Y(n747), 
	.B1(n805), 
	.B0(n210), 
	.A1(FE_OFN64_n258), 
	.A0(n804));
   OAI22X1 U478 (.Y(n748), 
	.B1(n804), 
	.B0(n210), 
	.A1(FE_OFN64_n258), 
	.A0(n803));
   OAI22X1 U479 (.Y(n749), 
	.B1(n803), 
	.B0(n210), 
	.A1(FE_OFN64_n258), 
	.A0(n802));
   OAI22X1 U480 (.Y(n750), 
	.B1(n802), 
	.B0(n210), 
	.A1(FE_PHN704_n258), 
	.A0(n801));
   OAI22X1 U481 (.Y(n751), 
	.B1(n801), 
	.B0(n210), 
	.A1(FE_PHN704_n258), 
	.A0(n800));
   OAI22X1 U482 (.Y(n752), 
	.B1(n800), 
	.B0(n210), 
	.A1(FE_PHN704_n258), 
	.A0(n799));
   OAI22X1 U483 (.Y(n753), 
	.B1(n799), 
	.B0(n210), 
	.A1(FE_PHN704_n258), 
	.A0(n798));
   OAI22X1 U484 (.Y(n754), 
	.B1(n798), 
	.B0(n210), 
	.A1(FE_PHN704_n258), 
	.A0(n797));
   OAI22X1 U485 (.Y(n755), 
	.B1(n797), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n796));
   OAI22X1 U486 (.Y(n756), 
	.B1(n796), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n795));
   OAI22X1 U487 (.Y(n757), 
	.B1(n795), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n794));
   OAI22X1 U488 (.Y(n758), 
	.B1(n794), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n793));
   OAI22X1 U489 (.Y(n759), 
	.B1(n793), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n792));
   OAI22X1 U490 (.Y(n760), 
	.B1(n792), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n791));
   OAI22X1 U491 (.Y(n761), 
	.B1(n791), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n790));
   OAI22X1 U492 (.Y(n762), 
	.B1(n790), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n789));
   OAI22X1 U493 (.Y(n763), 
	.B1(n789), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n788));
   OAI22X1 U494 (.Y(n764), 
	.B1(n788), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n787));
   OAI22X1 U495 (.Y(n765), 
	.B1(n787), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n786));
   OAI22X1 U496 (.Y(n766), 
	.B1(n786), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n785));
   OAI22X1 U497 (.Y(n767), 
	.B1(n785), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n784));
   OAI22X1 U498 (.Y(n768), 
	.B1(n784), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n783));
   OAI22X1 U499 (.Y(n769), 
	.B1(n783), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n782));
   OAI22X1 U500 (.Y(n770), 
	.B1(n782), 
	.B0(FE_OFN60_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n781));
   OAI22X1 U501 (.Y(n516), 
	.B1(n1036), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1035));
   OAI22X1 U502 (.Y(n548), 
	.B1(n1004), 
	.B0(FE_OFN63_n210), 
	.A1(FE_OFN65_n258), 
	.A0(n1003));
   OAI22X1 U503 (.Y(n580), 
	.B1(n972), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n971));
   OAI22X1 U504 (.Y(n612), 
	.B1(n940), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n939));
   OAI22X1 U505 (.Y(n644), 
	.B1(n908), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n907));
   OAI22X1 U506 (.Y(n676), 
	.B1(n876), 
	.B0(FE_OFN62_n210), 
	.A1(FE_OFN66_n258), 
	.A0(n875));
   OAI22X1 U507 (.Y(n708), 
	.B1(n844), 
	.B0(n210), 
	.A1(n52), 
	.A0(n843));
   OAI22X1 U508 (.Y(n740), 
	.B1(FE_PHN1243_n812), 
	.B0(FE_OFN61_n210), 
	.A1(FE_OFN64_n258), 
	.A0(n811));
   OAI2BB2X1 U517 (.Y(n547), 
	.B1(n1005), 
	.B0(FE_OFN62_n210), 
	.A1N(n171), 
	.A0N(plain_byte_in[0]));
   OAI2BB2X1 U518 (.Y(n579), 
	.B1(n973), 
	.B0(FE_OFN63_n210), 
	.A1N(FE_OFN63_n210), 
	.A0N(plain_byte_in[1]));
   OAI2BB2X1 U519 (.Y(n611), 
	.B1(n941), 
	.B0(FE_OFN63_n210), 
	.A1N(FE_OFN63_n210), 
	.A0N(plain_byte_in[2]));
   OAI2BB2X1 U520 (.Y(n643), 
	.B1(n909), 
	.B0(n210), 
	.A1N(n210), 
	.A0N(plain_byte_in[3]));
   OAI2BB2X1 U521 (.Y(n675), 
	.B1(n877), 
	.B0(n210), 
	.A1N(n210), 
	.A0N(plain_byte_in[4]));
   OAI2BB2X1 U522 (.Y(n707), 
	.B1(n845), 
	.B0(n210), 
	.A1N(n210), 
	.A0N(plain_byte_in[5]));
   OAI2BB2X1 U523 (.Y(n739), 
	.B1(n813), 
	.B0(n210), 
	.A1N(n210), 
	.A0N(plain_byte_in[6]));
   OAI2BB2X1 U524 (.Y(n771), 
	.B1(n781), 
	.B0(n210), 
	.A1N(n210), 
	.A0N(plain_byte_in[7]));
   NAND2BX1 U525 (.Y(n258), 
	.B(FE_PHN2804_pbv1), 
	.AN(FE_PHN2800_pbv0));
   NAND2BX2 U526 (.Y(n1), 
	.B(pf1), 
	.AN(FE_PHN2801_pf0));
   OAI2BB2X1 U527 (.Y(n260), 
	.B1(n1005), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[0]));
   OAI2BB2X1 U528 (.Y(n261), 
	.B1(n973), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[1]));
   OAI2BB2X1 U529 (.Y(n262), 
	.B1(n941), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[2]));
   OAI2BB2X1 U530 (.Y(n263), 
	.B1(n909), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[3]));
   OAI2BB2X1 U531 (.Y(n264), 
	.B1(n877), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[4]));
   OAI2BB2X1 U532 (.Y(n265), 
	.B1(n845), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[5]));
   OAI2BB2X1 U533 (.Y(n266), 
	.B1(n813), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[6]));
   OAI2BB2X1 U534 (.Y(n267), 
	.B1(n781), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[7]));
   OAI2BB2X1 U535 (.Y(n268), 
	.B1(n1006), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[8]));
   OAI2BB2X1 U536 (.Y(n269), 
	.B1(n974), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[9]));
   OAI2BB2X1 U537 (.Y(n270), 
	.B1(n942), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[10]));
   OAI2BB2X1 U538 (.Y(n271), 
	.B1(n910), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[11]));
   OAI2BB2X1 U539 (.Y(n272), 
	.B1(n878), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[12]));
   OAI2BB2X1 U540 (.Y(n273), 
	.B1(n846), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[13]));
   OAI2BB2X1 U541 (.Y(n274), 
	.B1(n814), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[14]));
   OAI2BB2X1 U542 (.Y(n275), 
	.B1(n782), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[15]));
   OAI2BB2X1 U543 (.Y(n276), 
	.B1(n1007), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[16]));
   OAI2BB2X1 U544 (.Y(n277), 
	.B1(n975), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[17]));
   OAI2BB2X1 U545 (.Y(n278), 
	.B1(n943), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[18]));
   OAI2BB2X1 U546 (.Y(n279), 
	.B1(n911), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[19]));
   OAI2BB2X1 U547 (.Y(n280), 
	.B1(n879), 
	.B0(FE_OFN71_n1), 
	.A1N(FE_OFN71_n1), 
	.A0N(plain_key_out[20]));
   OAI2BB2X1 U548 (.Y(n281), 
	.B1(n847), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[21]));
   OAI2BB2X1 U549 (.Y(n282), 
	.B1(n815), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[22]));
   OAI2BB2X1 U550 (.Y(n283), 
	.B1(n783), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[23]));
   OAI2BB2X1 U551 (.Y(n284), 
	.B1(n1008), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[24]));
   OAI2BB2X1 U552 (.Y(n285), 
	.B1(n976), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[25]));
   OAI2BB2X1 U553 (.Y(n286), 
	.B1(n944), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[26]));
   OAI2BB2X1 U554 (.Y(n287), 
	.B1(n912), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[27]));
   OAI2BB2X1 U555 (.Y(n288), 
	.B1(n880), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[28]));
   OAI2BB2X1 U556 (.Y(n289), 
	.B1(n848), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[29]));
   OAI2BB2X1 U557 (.Y(n290), 
	.B1(n816), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[30]));
   OAI2BB2X1 U558 (.Y(n291), 
	.B1(n784), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[31]));
   OAI2BB2X1 U559 (.Y(n292), 
	.B1(n1009), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[32]));
   OAI2BB2X1 U560 (.Y(n293), 
	.B1(n977), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[33]));
   OAI2BB2X1 U561 (.Y(n294), 
	.B1(n945), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[34]));
   OAI2BB2X1 U562 (.Y(n295), 
	.B1(n913), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[35]));
   OAI2BB2X1 U563 (.Y(n296), 
	.B1(n881), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[36]));
   OAI2BB2X1 U564 (.Y(n297), 
	.B1(n849), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[37]));
   OAI2BB2X1 U565 (.Y(n298), 
	.B1(n817), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[38]));
   OAI2BB2X1 U566 (.Y(n299), 
	.B1(n785), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[39]));
   OAI2BB2X1 U567 (.Y(n300), 
	.B1(n1010), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[40]));
   OAI2BB2X1 U568 (.Y(n301), 
	.B1(n978), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[41]));
   OAI2BB2X1 U569 (.Y(n302), 
	.B1(n946), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[42]));
   OAI2BB2X1 U570 (.Y(n303), 
	.B1(n914), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[43]));
   OAI2BB2X1 U571 (.Y(n304), 
	.B1(n882), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[44]));
   OAI2BB2X1 U572 (.Y(n305), 
	.B1(n850), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[45]));
   OAI2BB2X1 U573 (.Y(n306), 
	.B1(n818), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[46]));
   OAI2BB2X1 U574 (.Y(n307), 
	.B1(n786), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[47]));
   OAI2BB2X1 U575 (.Y(n308), 
	.B1(n1011), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[48]));
   OAI2BB2X1 U576 (.Y(n309), 
	.B1(n979), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[49]));
   OAI2BB2X1 U577 (.Y(n310), 
	.B1(n947), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[50]));
   OAI2BB2X1 U578 (.Y(n311), 
	.B1(n915), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[51]));
   OAI2BB2X1 U579 (.Y(n312), 
	.B1(n883), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[52]));
   OAI2BB2X1 U580 (.Y(n313), 
	.B1(n851), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[53]));
   OAI2BB2X1 U581 (.Y(n314), 
	.B1(n819), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[54]));
   OAI2BB2X1 U582 (.Y(n315), 
	.B1(n787), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[55]));
   OAI2BB2X1 U583 (.Y(n316), 
	.B1(n1012), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[56]));
   OAI2BB2X1 U584 (.Y(n317), 
	.B1(n980), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[57]));
   OAI2BB2X1 U585 (.Y(n318), 
	.B1(n948), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[58]));
   OAI2BB2X1 U586 (.Y(n319), 
	.B1(n916), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[59]));
   OAI2BB2X1 U587 (.Y(n320), 
	.B1(n884), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[60]));
   OAI2BB2X1 U588 (.Y(n321), 
	.B1(n852), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[61]));
   OAI2BB2X1 U589 (.Y(n322), 
	.B1(n820), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[62]));
   OAI2BB2X1 U590 (.Y(n323), 
	.B1(n788), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[63]));
   OAI2BB2X1 U591 (.Y(n324), 
	.B1(n1013), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[64]));
   OAI2BB2X1 U592 (.Y(n325), 
	.B1(n981), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[65]));
   OAI2BB2X1 U593 (.Y(n326), 
	.B1(n949), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[66]));
   OAI2BB2X1 U594 (.Y(n327), 
	.B1(n917), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[67]));
   OAI2BB2X1 U595 (.Y(n328), 
	.B1(n885), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[68]));
   OAI2BB2X1 U596 (.Y(n329), 
	.B1(n853), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[69]));
   OAI2BB2X1 U597 (.Y(n330), 
	.B1(n821), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[70]));
   OAI2BB2X1 U598 (.Y(n331), 
	.B1(n789), 
	.B0(FE_OFN71_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[71]));
   OAI2BB2X1 U599 (.Y(n332), 
	.B1(n1014), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[72]));
   OAI2BB2X1 U600 (.Y(n333), 
	.B1(n982), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[73]));
   OAI2BB2X1 U601 (.Y(n334), 
	.B1(n950), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[74]));
   OAI2BB2X1 U602 (.Y(n335), 
	.B1(n918), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[75]));
   OAI2BB2X1 U603 (.Y(n336), 
	.B1(n886), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[76]));
   OAI2BB2X1 U604 (.Y(n337), 
	.B1(n854), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[77]));
   OAI2BB2X1 U605 (.Y(n338), 
	.B1(n822), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[78]));
   OAI2BB2X1 U606 (.Y(n339), 
	.B1(n790), 
	.B0(FE_OFN71_n1), 
	.A1N(FE_OFN71_n1), 
	.A0N(plain_key_out[79]));
   OAI2BB2X1 U607 (.Y(n340), 
	.B1(n1015), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[80]));
   OAI2BB2X1 U608 (.Y(n341), 
	.B1(n983), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[81]));
   OAI2BB2X1 U609 (.Y(n342), 
	.B1(n951), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[82]));
   OAI2BB2X1 U610 (.Y(n343), 
	.B1(n919), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[83]));
   OAI2BB2X1 U611 (.Y(n344), 
	.B1(n887), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[84]));
   OAI2BB2X1 U612 (.Y(n345), 
	.B1(n855), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[85]));
   OAI2BB2X1 U613 (.Y(n346), 
	.B1(n823), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[86]));
   OAI2BB2X1 U614 (.Y(n347), 
	.B1(n791), 
	.B0(FE_OFN71_n1), 
	.A1N(FE_OFN71_n1), 
	.A0N(plain_key_out[87]));
   OAI2BB2X1 U615 (.Y(n348), 
	.B1(n1016), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[88]));
   OAI2BB2X1 U616 (.Y(n349), 
	.B1(n984), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[89]));
   OAI2BB2X1 U617 (.Y(n350), 
	.B1(n952), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[90]));
   OAI2BB2X1 U618 (.Y(n351), 
	.B1(n920), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[91]));
   OAI2BB2X1 U619 (.Y(n352), 
	.B1(n888), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[92]));
   OAI2BB2X1 U620 (.Y(n353), 
	.B1(n856), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[93]));
   OAI2BB2X1 U621 (.Y(n354), 
	.B1(n824), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[94]));
   OAI2BB2X1 U622 (.Y(n355), 
	.B1(n792), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[95]));
   OAI2BB2X1 U623 (.Y(n356), 
	.B1(n1017), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[96]));
   OAI2BB2X1 U624 (.Y(n357), 
	.B1(n985), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[97]));
   OAI2BB2X1 U625 (.Y(n358), 
	.B1(n953), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[98]));
   OAI2BB2X1 U626 (.Y(n359), 
	.B1(n921), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[99]));
   OAI2BB2X1 U627 (.Y(n360), 
	.B1(n889), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[100]));
   OAI2BB2X1 U628 (.Y(n361), 
	.B1(n857), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[101]));
   OAI2BB2X1 U629 (.Y(n362), 
	.B1(n825), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[102]));
   OAI2BB2X1 U630 (.Y(n363), 
	.B1(n793), 
	.B0(FE_OFN71_n1), 
	.A1N(FE_OFN71_n1), 
	.A0N(plain_key_out[103]));
   OAI2BB2X1 U631 (.Y(n364), 
	.B1(n1018), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[104]));
   OAI2BB2X1 U632 (.Y(n365), 
	.B1(n986), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[105]));
   OAI2BB2X1 U633 (.Y(n366), 
	.B1(n954), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[106]));
   OAI2BB2X1 U634 (.Y(n367), 
	.B1(n922), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[107]));
   OAI2BB2X1 U635 (.Y(n368), 
	.B1(n890), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[108]));
   OAI2BB2X1 U636 (.Y(n369), 
	.B1(n858), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[109]));
   OAI2BB2X1 U637 (.Y(n370), 
	.B1(n826), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[110]));
   OAI2BB2X1 U638 (.Y(n371), 
	.B1(n794), 
	.B0(FE_OFN71_n1), 
	.A1N(FE_OFN71_n1), 
	.A0N(plain_key_out[111]));
   OAI2BB2X1 U639 (.Y(n372), 
	.B1(n1019), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[112]));
   OAI2BB2X1 U640 (.Y(n373), 
	.B1(n987), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[113]));
   OAI2BB2X1 U641 (.Y(n374), 
	.B1(n955), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[114]));
   OAI2BB2X1 U642 (.Y(n375), 
	.B1(n923), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[115]));
   OAI2BB2X1 U643 (.Y(n376), 
	.B1(n891), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[116]));
   OAI2BB2X1 U644 (.Y(n377), 
	.B1(n859), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[117]));
   OAI2BB2X1 U645 (.Y(n378), 
	.B1(n827), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[118]));
   OAI2BB2X1 U646 (.Y(n379), 
	.B1(n795), 
	.B0(FE_OFN71_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[119]));
   OAI2BB2X1 U647 (.Y(n380), 
	.B1(n1020), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[120]));
   OAI2BB2X1 U648 (.Y(n381), 
	.B1(n988), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[121]));
   OAI2BB2X1 U649 (.Y(n382), 
	.B1(n956), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[122]));
   OAI2BB2X1 U650 (.Y(n383), 
	.B1(n924), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[123]));
   OAI2BB2X1 U651 (.Y(n384), 
	.B1(n892), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[124]));
   OAI2BB2X1 U652 (.Y(n385), 
	.B1(n860), 
	.B0(FE_OFN70_n1), 
	.A1N(FE_OFN70_n1), 
	.A0N(plain_key_out[125]));
   OAI2BB2X1 U653 (.Y(n386), 
	.B1(n828), 
	.B0(FE_OFN68_n1), 
	.A1N(FE_OFN68_n1), 
	.A0N(plain_key_out[126]));
   OAI2BB2X1 U654 (.Y(n387), 
	.B1(n796), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[127]));
   OAI2BB2X1 U655 (.Y(n388), 
	.B1(n1021), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[128]));
   OAI2BB2X1 U656 (.Y(n389), 
	.B1(n989), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[129]));
   OAI2BB2X1 U657 (.Y(n390), 
	.B1(n957), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[130]));
   OAI2BB2X1 U658 (.Y(n391), 
	.B1(n925), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[131]));
   OAI2BB2X1 U659 (.Y(n392), 
	.B1(n893), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[132]));
   OAI2BB2X1 U660 (.Y(n393), 
	.B1(n861), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[133]));
   OAI2BB2X1 U661 (.Y(n394), 
	.B1(n829), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[134]));
   OAI2BB2X1 U662 (.Y(n395), 
	.B1(n797), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[135]));
   OAI2BB2X1 U663 (.Y(n396), 
	.B1(n1022), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[136]));
   OAI2BB2X1 U664 (.Y(n397), 
	.B1(n990), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[137]));
   OAI2BB2X1 U665 (.Y(n398), 
	.B1(n958), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[138]));
   OAI2BB2X1 U666 (.Y(n399), 
	.B1(n926), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[139]));
   OAI2BB2X1 U667 (.Y(n400), 
	.B1(n894), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[140]));
   OAI2BB2X1 U668 (.Y(n401), 
	.B1(n862), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[141]));
   OAI2BB2X1 U669 (.Y(n402), 
	.B1(n830), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[142]));
   OAI2BB2X1 U670 (.Y(n403), 
	.B1(n798), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[143]));
   OAI2BB2X1 U671 (.Y(n404), 
	.B1(n1023), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[144]));
   OAI2BB2X1 U672 (.Y(n405), 
	.B1(n991), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[145]));
   OAI2BB2X1 U673 (.Y(n406), 
	.B1(n959), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[146]));
   OAI2BB2X1 U674 (.Y(n407), 
	.B1(n927), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[147]));
   OAI2BB2X1 U675 (.Y(n408), 
	.B1(n895), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[148]));
   OAI2BB2X1 U676 (.Y(n409), 
	.B1(n863), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[149]));
   OAI2BB2X1 U677 (.Y(n410), 
	.B1(n831), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[150]));
   OAI2BB2X1 U678 (.Y(n411), 
	.B1(n799), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[151]));
   OAI2BB2X1 U679 (.Y(n412), 
	.B1(n1024), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[152]));
   OAI2BB2X1 U680 (.Y(n413), 
	.B1(n992), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[153]));
   OAI2BB2X1 U681 (.Y(n414), 
	.B1(n960), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[154]));
   OAI2BB2X1 U682 (.Y(n415), 
	.B1(n928), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[155]));
   OAI2BB2X1 U683 (.Y(n416), 
	.B1(n896), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[156]));
   OAI2BB2X1 U684 (.Y(n417), 
	.B1(n864), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[157]));
   OAI2BB2X1 U685 (.Y(n418), 
	.B1(n832), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[158]));
   OAI2BB2X1 U686 (.Y(n419), 
	.B1(n800), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[159]));
   OAI2BB2X1 U687 (.Y(n420), 
	.B1(n1025), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[160]));
   OAI2BB2X1 U688 (.Y(n421), 
	.B1(n993), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[161]));
   OAI2BB2X1 U689 (.Y(n422), 
	.B1(n961), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[162]));
   OAI2BB2X1 U690 (.Y(n423), 
	.B1(n929), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[163]));
   OAI2BB2X1 U691 (.Y(n424), 
	.B1(n897), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[164]));
   OAI2BB2X1 U692 (.Y(n425), 
	.B1(n865), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[165]));
   OAI2BB2X1 U693 (.Y(n426), 
	.B1(n833), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[166]));
   OAI2BB2X1 U694 (.Y(n427), 
	.B1(n801), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[167]));
   OAI2BB2X1 U695 (.Y(n428), 
	.B1(n1026), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[168]));
   OAI2BB2X1 U696 (.Y(n429), 
	.B1(n994), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[169]));
   OAI2BB2X1 U697 (.Y(n430), 
	.B1(n962), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[170]));
   OAI2BB2X1 U698 (.Y(n431), 
	.B1(n930), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[171]));
   OAI2BB2X1 U699 (.Y(n432), 
	.B1(n898), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[172]));
   OAI2BB2X1 U700 (.Y(n433), 
	.B1(n866), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[173]));
   OAI2BB2X1 U701 (.Y(n434), 
	.B1(n834), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[174]));
   OAI2BB2X1 U702 (.Y(n435), 
	.B1(n802), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[175]));
   OAI2BB2X1 U703 (.Y(n436), 
	.B1(n1027), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[176]));
   OAI2BB2X1 U704 (.Y(n437), 
	.B1(n995), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[177]));
   OAI2BB2X1 U705 (.Y(n438), 
	.B1(n963), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[178]));
   OAI2BB2X1 U706 (.Y(n439), 
	.B1(n931), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[179]));
   OAI2BB2X1 U707 (.Y(n440), 
	.B1(n899), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[180]));
   OAI2BB2X1 U708 (.Y(n441), 
	.B1(n867), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[181]));
   OAI2BB2X1 U709 (.Y(n442), 
	.B1(n835), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[182]));
   OAI2BB2X1 U710 (.Y(n443), 
	.B1(n803), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[183]));
   OAI2BB2X1 U711 (.Y(n444), 
	.B1(n1028), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[184]));
   OAI2BB2X1 U712 (.Y(n445), 
	.B1(n996), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[185]));
   OAI2BB2X1 U713 (.Y(n446), 
	.B1(n964), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[186]));
   OAI2BB2X1 U714 (.Y(n447), 
	.B1(n932), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[187]));
   OAI2BB2X1 U715 (.Y(n448), 
	.B1(n900), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[188]));
   OAI2BB2X1 U716 (.Y(n449), 
	.B1(n868), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[189]));
   OAI2BB2X1 U717 (.Y(n450), 
	.B1(n836), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[190]));
   OAI2BB2X1 U718 (.Y(n451), 
	.B1(n804), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[191]));
   OAI2BB2X1 U719 (.Y(n452), 
	.B1(n1029), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[192]));
   OAI2BB2X1 U720 (.Y(n453), 
	.B1(n997), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[193]));
   OAI2BB2X1 U721 (.Y(n454), 
	.B1(n965), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[194]));
   OAI2BB2X1 U722 (.Y(n455), 
	.B1(n933), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[195]));
   OAI2BB2X1 U723 (.Y(n456), 
	.B1(n901), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[196]));
   OAI2BB2X1 U724 (.Y(n457), 
	.B1(n869), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[197]));
   OAI2BB2X1 U725 (.Y(n458), 
	.B1(n837), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[198]));
   OAI2BB2X1 U726 (.Y(n459), 
	.B1(n805), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[199]));
   OAI2BB2X1 U727 (.Y(n460), 
	.B1(n1030), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[200]));
   OAI2BB2X1 U728 (.Y(n461), 
	.B1(n998), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[201]));
   OAI2BB2X1 U729 (.Y(n462), 
	.B1(n966), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[202]));
   OAI2BB2X1 U730 (.Y(n463), 
	.B1(n934), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[203]));
   OAI2BB2X1 U731 (.Y(n464), 
	.B1(n902), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[204]));
   OAI2BB2X1 U732 (.Y(n465), 
	.B1(n870), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[205]));
   OAI2BB2X1 U733 (.Y(n466), 
	.B1(n838), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[206]));
   OAI2BB2X1 U734 (.Y(n467), 
	.B1(n806), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[207]));
   OAI2BB2X1 U735 (.Y(n468), 
	.B1(n1031), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[208]));
   OAI2BB2X1 U736 (.Y(n469), 
	.B1(n999), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[209]));
   OAI2BB2X1 U737 (.Y(n470), 
	.B1(n967), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[210]));
   OAI2BB2X1 U738 (.Y(n471), 
	.B1(n935), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[211]));
   OAI2BB2X1 U739 (.Y(n472), 
	.B1(n903), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[212]));
   OAI2BB2X1 U740 (.Y(n473), 
	.B1(n871), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[213]));
   OAI2BB2X1 U741 (.Y(n474), 
	.B1(n839), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[214]));
   OAI2BB2X1 U742 (.Y(n475), 
	.B1(n807), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[215]));
   OAI2BB2X1 U743 (.Y(n476), 
	.B1(n1032), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[216]));
   OAI2BB2X1 U744 (.Y(n477), 
	.B1(n1000), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[217]));
   OAI2BB2X1 U745 (.Y(n478), 
	.B1(n968), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[218]));
   OAI2BB2X1 U746 (.Y(n479), 
	.B1(n936), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[219]));
   OAI2BB2X1 U747 (.Y(n480), 
	.B1(n904), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[220]));
   OAI2BB2X1 U748 (.Y(n481), 
	.B1(n872), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[221]));
   OAI2BB2X1 U749 (.Y(n482), 
	.B1(n840), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[222]));
   OAI2BB2X1 U750 (.Y(n483), 
	.B1(n808), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[223]));
   OAI2BB2X1 U751 (.Y(n484), 
	.B1(n1033), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[224]));
   OAI2BB2X1 U752 (.Y(n485), 
	.B1(n1001), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[225]));
   OAI2BB2X1 U753 (.Y(n486), 
	.B1(n969), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[226]));
   OAI2BB2X1 U754 (.Y(n487), 
	.B1(n937), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[227]));
   OAI2BB2X1 U755 (.Y(n488), 
	.B1(n905), 
	.B0(FE_OFN74_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[228]));
   OAI2BB2X1 U756 (.Y(n489), 
	.B1(n873), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[229]));
   OAI2BB2X1 U757 (.Y(n490), 
	.B1(n841), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[230]));
   OAI2BB2X1 U758 (.Y(n491), 
	.B1(n809), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[231]));
   OAI2BB2X1 U759 (.Y(n492), 
	.B1(n1034), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[232]));
   OAI2BB2X1 U760 (.Y(n493), 
	.B1(n1002), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[233]));
   OAI2BB2X1 U761 (.Y(n494), 
	.B1(n970), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[234]));
   OAI2BB2X1 U762 (.Y(n495), 
	.B1(n938), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN74_n1), 
	.A0N(plain_key_out[235]));
   OAI2BB2X1 U763 (.Y(n496), 
	.B1(n906), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[236]));
   OAI2BB2X1 U764 (.Y(n497), 
	.B1(n874), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[237]));
   OAI2BB2X1 U765 (.Y(n498), 
	.B1(n842), 
	.B0(FE_PHN119_n1), 
	.A1N(FE_PHN119_n1), 
	.A0N(plain_key_out[238]));
   OAI2BB2X1 U766 (.Y(n499), 
	.B1(n810), 
	.B0(FE_OFN71_n1), 
	.A1N(FE_OFN71_n1), 
	.A0N(plain_key_out[239]));
   OAI2BB2X1 U767 (.Y(n500), 
	.B1(n1035), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[240]));
   OAI2BB2X1 U768 (.Y(n501), 
	.B1(n1003), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[241]));
   OAI2BB2X1 U769 (.Y(n502), 
	.B1(n971), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[242]));
   OAI2BB2X1 U770 (.Y(n503), 
	.B1(n939), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[243]));
   OAI2BB2X1 U771 (.Y(n504), 
	.B1(n907), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[244]));
   OAI2BB2X1 U772 (.Y(n505), 
	.B1(n875), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[245]));
   OAI2BB2X1 U773 (.Y(n506), 
	.B1(n843), 
	.B0(FE_OFN71_n1), 
	.A1N(FE_OFN71_n1), 
	.A0N(plain_key_out[246]));
   OAI2BB2X1 U774 (.Y(n507), 
	.B1(n811), 
	.B0(FE_OFN71_n1), 
	.A1N(FE_OFN71_n1), 
	.A0N(plain_key_out[247]));
   OAI2BB2X1 U775 (.Y(n508), 
	.B1(n1036), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[248]));
   OAI2BB2X1 U776 (.Y(n509), 
	.B1(n1004), 
	.B0(FE_OFN75_n1), 
	.A1N(FE_OFN75_n1), 
	.A0N(plain_key_out[249]));
   OAI2BB2X1 U777 (.Y(n510), 
	.B1(n972), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[250]));
   OAI2BB2X1 U778 (.Y(n511), 
	.B1(n940), 
	.B0(FE_OFN72_n1), 
	.A1N(FE_OFN72_n1), 
	.A0N(plain_key_out[251]));
   OAI2BB2X1 U779 (.Y(n512), 
	.B1(n908), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[252]));
   OAI2BB2X1 U780 (.Y(n513), 
	.B1(n876), 
	.B0(FE_OFN73_n1), 
	.A1N(FE_OFN73_n1), 
	.A0N(plain_key_out[253]));
   OAI2BB2X1 U781 (.Y(n514), 
	.B1(n844), 
	.B0(FE_OFN69_n1), 
	.A1N(FE_OFN69_n1), 
	.A0N(plain_key_out[254]));
   OAI2BB2X1 U782 (.Y(n515), 
	.B1(FE_PHN1243_n812), 
	.B0(FE_OFN71_n1), 
	.A1N(FE_OFN71_n1), 
	.A0N(plain_key_out[255]));
   INVX1 U783 (.Y(n1005), 
	.A(FE_PHN3391_plain_text_0_));
   INVX1 U784 (.Y(n973), 
	.A(FE_PHN1462_plain_text_1_));
   INVX1 U785 (.Y(n941), 
	.A(FE_PHN1460_plain_text_2_));
   INVX1 U786 (.Y(n909), 
	.A(FE_PHN1210_plain_text_3_));
   INVX1 U787 (.Y(n877), 
	.A(FE_PHN2888_plain_text_4_));
   INVX1 U788 (.Y(n845), 
	.A(FE_PHN3079_plain_text_5_));
   INVX1 U789 (.Y(n813), 
	.A(FE_PHN1450_plain_text_6_));
   INVX1 U790 (.Y(n781), 
	.A(FE_PHN3171_plain_text_7_));
   INVX1 U791 (.Y(n1035), 
	.A(FE_PHN1400_plain_text_240_));
   INVX1 U792 (.Y(n1034), 
	.A(FE_PHN2031_plain_text_232_));
   INVX1 U793 (.Y(n1033), 
	.A(FE_PHN1368_plain_text_224_));
   INVX1 U794 (.Y(n1032), 
	.A(FE_PHN3136_plain_text_216_));
   INVX1 U795 (.Y(n1031), 
	.A(FE_PHN3008_plain_text_208_));
   INVX1 U796 (.Y(n1030), 
	.A(FE_PHN3040_plain_text_200_));
   INVX1 U797 (.Y(n1029), 
	.A(FE_PHN1108_plain_text_192_));
   INVX1 U798 (.Y(n1028), 
	.A(FE_PHN2027_plain_text_184_));
   INVX1 U799 (.Y(n1027), 
	.A(FE_PHN1350_plain_text_176_));
   INVX1 U800 (.Y(n1026), 
	.A(FE_PHN1163_plain_text_168_));
   INVX1 U801 (.Y(n1025), 
	.A(FE_PHN2019_plain_text_160_));
   INVX1 U802 (.Y(n1024), 
	.A(FE_PHN1194_plain_text_152_));
   INVX1 U803 (.Y(n1023), 
	.A(FE_PHN2025_plain_text_144_));
   INVX1 U804 (.Y(n1022), 
	.A(FE_PHN1364_plain_text_136_));
   INVX1 U805 (.Y(n1021), 
	.A(FE_PHN3121_plain_text_128_));
   INVX1 U806 (.Y(n1020), 
	.A(FE_PHN1148_plain_text_120_));
   INVX1 U807 (.Y(n1019), 
	.A(FE_PHN3030_plain_text_112_));
   INVX1 U808 (.Y(n1018), 
	.A(FE_PHN1112_plain_text_104_));
   INVX1 U809 (.Y(n1017), 
	.A(FE_PHN2973_plain_text_96_));
   INVX1 U810 (.Y(n1016), 
	.A(FE_PHN2958_plain_text_88_));
   INVX1 U811 (.Y(n1015), 
	.A(FE_PHN2977_plain_text_80_));
   INVX1 U812 (.Y(n1014), 
	.A(FE_PHN3124_plain_text_72_));
   INVX1 U813 (.Y(n1013), 
	.A(FE_PHN2861_plain_text_64_));
   INVX1 U814 (.Y(n1012), 
	.A(FE_PHN1122_plain_text_56_));
   INVX1 U815 (.Y(n1011), 
	.A(FE_PHN1382_plain_text_48_));
   INVX1 U816 (.Y(n1010), 
	.A(FE_PHN2884_plain_text_40_));
   INVX1 U817 (.Y(n1009), 
	.A(FE_PHN1355_plain_text_32_));
   INVX1 U818 (.Y(n1008), 
	.A(FE_PHN3054_plain_text_24_));
   INVX1 U819 (.Y(n1007), 
	.A(FE_PHN2880_plain_text_16_));
   INVX1 U820 (.Y(n1006), 
	.A(FE_PHN1201_plain_text_8_));
   INVX1 U821 (.Y(n1003), 
	.A(FE_PHN1147_plain_text_241_));
   INVX1 U822 (.Y(n1002), 
	.A(FE_PHN2012_plain_text_233_));
   INVX1 U823 (.Y(n1001), 
	.A(FE_PHN3355_plain_text_225_));
   INVX1 U824 (.Y(n1000), 
	.A(FE_PHN1099_plain_text_217_));
   INVX1 U825 (.Y(n999), 
	.A(FE_PHN2026_plain_text_209_));
   INVX1 U826 (.Y(n998), 
	.A(FE_PHN1329_plain_text_201_));
   INVX1 U827 (.Y(n997), 
	.A(FE_PHN3311_plain_text_193_));
   INVX1 U828 (.Y(n996), 
	.A(FE_PHN2023_plain_text_185_));
   INVX1 U829 (.Y(n995), 
	.A(FE_PHN1385_plain_text_177_));
   INVX1 U830 (.Y(n994), 
	.A(FE_PHN3131_plain_text_169_));
   INVX1 U831 (.Y(n993), 
	.A(FE_PHN1127_plain_text_161_));
   INVX1 U832 (.Y(n992), 
	.A(FE_PHN2029_plain_text_153_));
   INVX1 U833 (.Y(n991), 
	.A(FE_PHN1396_plain_text_145_));
   INVX1 U834 (.Y(n990), 
	.A(FE_PHN1325_plain_text_137_));
   INVX1 U835 (.Y(n989), 
	.A(FE_PHN3112_plain_text_129_));
   INVX1 U836 (.Y(n988), 
	.A(FE_PHN5234_plain_text_121_));
   INVX1 U837 (.Y(n987), 
	.A(FE_PHN2945_plain_text_113_));
   INVX1 U838 (.Y(n986), 
	.A(FE_PHN1078_plain_text_105_));
   INVX1 U839 (.Y(n985), 
	.A(FE_PHN2952_plain_text_97_));
   INVX1 U840 (.Y(n984), 
	.A(FE_PHN1142_plain_text_89_));
   INVX1 U841 (.Y(n983), 
	.A(FE_PHN1343_plain_text_81_));
   INVX1 U842 (.Y(n982), 
	.A(FE_PHN1344_plain_text_73_));
   INVX1 U843 (.Y(n981), 
	.A(FE_PHN1369_plain_text_65_));
   INVX1 U844 (.Y(n980), 
	.A(FE_PHN1111_plain_text_57_));
   INVX1 U845 (.Y(n979), 
	.A(FE_PHN1089_plain_text_49_));
   INVX1 U846 (.Y(n978), 
	.A(FE_PHN2017_plain_text_41_));
   INVX1 U847 (.Y(n977), 
	.A(FE_PHN1082_plain_text_33_));
   INVX1 U848 (.Y(n976), 
	.A(FE_PHN3165_plain_text_25_));
   INVX1 U849 (.Y(n975), 
	.A(FE_PHN3044_plain_text_17_));
   INVX1 U850 (.Y(n974), 
	.A(FE_PHN2971_plain_text_9_));
   INVX1 U851 (.Y(n971), 
	.A(FE_PHN2020_plain_text_242_));
   INVX1 U852 (.Y(n970), 
	.A(FE_PHN3096_plain_text_234_));
   INVX1 U853 (.Y(n969), 
	.A(FE_PHN2032_plain_text_226_));
   INVX1 U854 (.Y(n968), 
	.A(FE_PHN1389_plain_text_218_));
   INVX1 U855 (.Y(n967), 
	.A(FE_PHN3152_plain_text_210_));
   INVX1 U856 (.Y(n966), 
	.A(FE_PHN3031_plain_text_202_));
   INVX1 U857 (.Y(n965), 
	.A(FE_PHN3012_plain_text_194_));
   INVX1 U858 (.Y(n964), 
	.A(FE_PHN2994_plain_text_186_));
   INVX1 U859 (.Y(n963), 
	.A(FE_PHN3148_plain_text_178_));
   INVX1 U860 (.Y(n962), 
	.A(FE_PHN1365_plain_text_170_));
   INVX1 U861 (.Y(n961), 
	.A(FE_PHN3099_plain_text_162_));
   INVX1 U862 (.Y(n960), 
	.A(FE_PHN2034_plain_text_154_));
   INVX1 U863 (.Y(n959), 
	.A(FE_PHN3369_plain_text_146_));
   INVX1 U864 (.Y(n958), 
	.A(FE_PHN3137_plain_text_138_));
   INVX1 U865 (.Y(n957), 
	.A(FE_PHN1124_plain_text_130_));
   INVX1 U866 (.Y(n956), 
	.A(FE_PHN1438_plain_text_122_));
   INVX1 U867 (.Y(n955), 
	.A(FE_PHN3052_plain_text_114_));
   INVX1 U868 (.Y(n954), 
	.A(FE_PHN2991_plain_text_106_));
   INVX1 U869 (.Y(n953), 
	.A(FE_PHN2992_plain_text_98_));
   INVX1 U870 (.Y(n952), 
	.A(FE_PHN3017_plain_text_90_));
   INVX1 U871 (.Y(n951), 
	.A(FE_PHN1097_plain_text_82_));
   INVX1 U872 (.Y(n950), 
	.A(FE_PHN1342_plain_text_74_));
   INVX1 U873 (.Y(n949), 
	.A(FE_PHN1114_plain_text_66_));
   INVX1 U874 (.Y(n948), 
	.A(FE_PHN1384_plain_text_58_));
   INVX1 U875 (.Y(n947), 
	.A(FE_PHN2867_plain_text_50_));
   INVX1 U876 (.Y(n946), 
	.A(FE_PHN1359_plain_text_42_));
   INVX1 U877 (.Y(n945), 
	.A(FE_PHN2932_plain_text_34_));
   INVX1 U878 (.Y(n944), 
	.A(FE_PHN2874_plain_text_26_));
   INVX1 U879 (.Y(n943), 
	.A(FE_PHN3382_plain_text_18_));
   INVX1 U880 (.Y(n942), 
	.A(FE_PHN3103_plain_text_10_));
   INVX1 U881 (.Y(n939), 
	.A(FE_PHN3336_plain_text_243_));
   INVX1 U882 (.Y(n938), 
	.A(FE_PHN2035_plain_text_235_));
   INVX1 U883 (.Y(n937), 
	.A(FE_PHN3101_plain_text_227_));
   INVX1 U884 (.Y(n936), 
	.A(FE_PHN2030_plain_text_219_));
   INVX1 U885 (.Y(n935), 
	.A(FE_PHN1118_plain_text_211_));
   INVX1 U886 (.Y(n934), 
	.A(FE_PHN1180_plain_text_203_));
   INVX1 U887 (.Y(n933), 
	.A(FE_PHN2014_plain_text_195_));
   INVX1 U888 (.Y(n932), 
	.A(FE_PHN1417_plain_text_187_));
   INVX1 U889 (.Y(n931), 
	.A(FE_PHN1430_plain_text_179_));
   INVX1 U890 (.Y(n930), 
	.A(FE_PHN1411_plain_text_171_));
   INVX1 U891 (.Y(n929), 
	.A(FE_PHN3363_plain_text_163_));
   INVX1 U892 (.Y(n928), 
	.A(FE_PHN882_plain_text_155_));
   INVX1 U893 (.Y(n927), 
	.A(FE_PHN1427_plain_text_147_));
   INVX1 U894 (.Y(n926), 
	.A(FE_PHN3576_plain_text_139_));
   INVX1 U895 (.Y(n925), 
	.A(FE_PHN3025_plain_text_131_));
   INVX1 U896 (.Y(n924), 
	.A(FE_PHN1452_plain_text_123_));
   INVX1 U897 (.Y(n923), 
	.A(FE_PHN1145_plain_text_115_));
   INVX1 U898 (.Y(n922), 
	.A(FE_PHN3037_plain_text_107_));
   INVX1 U899 (.Y(n921), 
	.A(FE_PHN3020_plain_text_99_));
   INVX1 U900 (.Y(n920), 
	.A(FE_PHN3015_plain_text_91_));
   INVX1 U901 (.Y(n919), 
	.A(FE_PHN2965_plain_text_83_));
   INVX1 U902 (.Y(n918), 
	.A(FE_PHN3092_plain_text_75_));
   INVX1 U903 (.Y(n917), 
	.A(FE_PHN2015_plain_text_67_));
   INVX1 U904 (.Y(n916), 
	.A(FE_PHN3376_plain_text_59_));
   INVX1 U905 (.Y(n915), 
	.A(FE_PHN2929_plain_text_51_));
   INVX1 U906 (.Y(n914), 
	.A(FE_PHN864_plain_text_43_));
   INVX1 U907 (.Y(n913), 
	.A(FE_PHN2016_plain_text_35_));
   INVX1 U908 (.Y(n912), 
	.A(FE_PHN1091_plain_text_27_));
   INVX1 U909 (.Y(n911), 
	.A(FE_PHN2871_plain_text_19_));
   INVX1 U910 (.Y(n910), 
	.A(FE_PHN1170_plain_text_11_));
   INVX1 U911 (.Y(n907), 
	.A(FE_PHN1331_plain_text_244_));
   INVX1 U912 (.Y(n906), 
	.A(FE_PHN2953_plain_text_236_));
   INVX1 U913 (.Y(n905), 
	.A(FE_PHN1398_plain_text_228_));
   INVX1 U914 (.Y(n904), 
	.A(FE_PHN1105_plain_text_220_));
   INVX1 U915 (.Y(n903), 
	.A(FE_PHN860_plain_text_212_));
   INVX1 U916 (.Y(n902), 
	.A(FE_PHN3588_plain_text_204_));
   INVX1 U917 (.Y(n901), 
	.A(FE_PHN3367_plain_text_196_));
   INVX1 U918 (.Y(n900), 
	.A(FE_PHN1059_plain_text_188_));
   INVX1 U919 (.Y(n899), 
	.A(FE_PHN830_plain_text_180_));
   INVX1 U920 (.Y(n898), 
	.A(FE_PHN2028_plain_text_172_));
   INVX1 U921 (.Y(n897), 
	.A(FE_PHN1102_plain_text_164_));
   INVX1 U922 (.Y(n896), 
	.A(FE_PHN1160_plain_text_156_));
   INVX1 U923 (.Y(n895), 
	.A(FE_PHN2964_plain_text_148_));
   INVX1 U924 (.Y(n894), 
	.A(FE_PHN2868_plain_text_140_));
   INVX1 U925 (.Y(n893), 
	.A(FE_PHN1440_plain_text_132_));
   INVX1 U926 (.Y(n892), 
	.A(FE_PHN2037_plain_text_124_));
   INVX1 U927 (.Y(n891), 
	.A(FE_PHN1206_plain_text_116_));
   INVX1 U928 (.Y(n890), 
	.A(FE_PHN1120_plain_text_108_));
   INVX1 U929 (.Y(n889), 
	.A(FE_PHN2942_plain_text_100_));
   INVX1 U930 (.Y(n888), 
	.A(FE_PHN2998_plain_text_92_));
   INVX1 U931 (.Y(n887), 
	.A(FE_PHN1119_plain_text_84_));
   INVX1 U932 (.Y(n886), 
	.A(FE_PHN1103_plain_text_76_));
   INVX1 U933 (.Y(n885), 
	.A(FE_PHN1320_plain_text_68_));
   INVX1 U934 (.Y(n884), 
	.A(FE_PHN1176_plain_text_60_));
   INVX1 U935 (.Y(n883), 
	.A(FE_PHN1073_plain_text_52_));
   INVX1 U936 (.Y(n882), 
	.A(FE_PHN2950_plain_text_44_));
   INVX1 U937 (.Y(n881), 
	.A(FE_PHN2875_plain_text_36_));
   INVX1 U938 (.Y(n880), 
	.A(FE_PHN5257_plain_text_28_));
   INVX1 U939 (.Y(n879), 
	.A(FE_PHN2860_plain_text_20_));
   INVX1 U940 (.Y(n878), 
	.A(FE_PHN5242_plain_text_12_));
   INVX1 U941 (.Y(n875), 
	.A(FE_PHN2010_plain_text_245_));
   INVX1 U942 (.Y(n874), 
	.A(FE_PHN835_plain_text_237_));
   INVX1 U943 (.Y(n873), 
	.A(FE_PHN2021_plain_text_229_));
   INVX1 U944 (.Y(n872), 
	.A(FE_PHN1130_plain_text_221_));
   INVX1 U945 (.Y(n871), 
	.A(FE_PHN2969_plain_text_213_));
   INVX1 U946 (.Y(n870), 
	.A(FE_PHN3153_plain_text_205_));
   INVX1 U947 (.Y(n869), 
	.A(FE_PHN2857_plain_text_197_));
   INVX1 U948 (.Y(n868), 
	.A(FE_PHN3154_plain_text_189_));
   INVX1 U949 (.Y(n867), 
	.A(FE_PHN1169_plain_text_181_));
   INVX1 U950 (.Y(n866), 
	.A(FE_PHN1168_plain_text_173_));
   INVX1 U951 (.Y(n865), 
	.A(FE_PHN2024_plain_text_165_));
   INVX1 U952 (.Y(n864), 
	.A(FE_PHN3389_plain_text_157_));
   INVX1 U953 (.Y(n863), 
	.A(FE_PHN3010_plain_text_149_));
   INVX1 U954 (.Y(n862), 
	.A(FE_PHN1327_plain_text_141_));
   INVX1 U955 (.Y(n861), 
	.A(FE_PHN3386_plain_text_133_));
   INVX1 U956 (.Y(n860), 
	.A(FE_PHN5072_plain_text_125_));
   INVX1 U957 (.Y(n859), 
	.A(FE_PHN1173_plain_text_117_));
   INVX1 U958 (.Y(n858), 
	.A(FE_PHN3043_plain_text_109_));
   INVX1 U959 (.Y(n857), 
	.A(FE_PHN3038_plain_text_101_));
   INVX1 U960 (.Y(n856), 
	.A(FE_PHN1167_plain_text_93_));
   INVX1 U961 (.Y(n855), 
	.A(FE_PHN2995_plain_text_85_));
   INVX1 U962 (.Y(n854), 
	.A(FE_PHN2882_plain_text_77_));
   INVX1 U963 (.Y(n853), 
	.A(FE_PHN3164_plain_text_69_));
   INVX1 U964 (.Y(n852), 
	.A(FE_PHN1187_plain_text_61_));
   INVX1 U965 (.Y(n851), 
	.A(FE_PHN2926_plain_text_53_));
   INVX1 U966 (.Y(n850), 
	.A(FE_PHN1149_plain_text_45_));
   INVX1 U967 (.Y(n849), 
	.A(FE_PHN2978_plain_text_37_));
   INVX1 U968 (.Y(n848), 
	.A(FE_PHN3034_plain_text_29_));
   INVX1 U969 (.Y(n847), 
	.A(FE_PHN1133_plain_text_21_));
   INVX1 U970 (.Y(n846), 
	.A(FE_PHN2876_plain_text_13_));
   INVX1 U971 (.Y(n843), 
	.A(FE_PHN3065_plain_text_246_));
   INVX1 U972 (.Y(n842), 
	.A(FE_PHN2033_plain_text_238_));
   INVX1 U973 (.Y(n841), 
	.A(FE_PHN1346_plain_text_230_));
   INVX1 U974 (.Y(n840), 
	.A(FE_PHN2966_plain_text_222_));
   INVX1 U975 (.Y(n839), 
	.A(FE_PHN1447_plain_text_214_));
   INVX1 U976 (.Y(n838), 
	.A(FE_PHN3143_plain_text_206_));
   INVX1 U977 (.Y(n837), 
	.A(FE_PHN1358_plain_text_198_));
   INVX1 U978 (.Y(n836), 
	.A(FE_PHN3045_plain_text_190_));
   INVX1 U979 (.Y(n835), 
	.A(FE_PHN3169_plain_text_182_));
   INVX1 U980 (.Y(n834), 
	.A(FE_PHN1403_plain_text_174_));
   INVX1 U981 (.Y(n833), 
	.A(FE_PHN1039_plain_text_166_));
   INVX1 U982 (.Y(n832), 
	.A(FE_PHN1152_plain_text_158_));
   INVX1 U983 (.Y(n831), 
	.A(FE_PHN3097_plain_text_150_));
   INVX1 U984 (.Y(n830), 
	.A(FE_PHN1341_plain_text_142_));
   INVX1 U985 (.Y(n829), 
	.A(FE_PHN2877_plain_text_134_));
   INVX1 U986 (.Y(n828), 
	.A(FE_PHN1436_plain_text_126_));
   INVX1 U987 (.Y(n827), 
	.A(FE_PHN3102_plain_text_118_));
   INVX1 U988 (.Y(n826), 
	.A(FE_PHN1123_plain_text_110_));
   INVX1 U989 (.Y(n825), 
	.A(FE_PHN2981_plain_text_102_));
   INVX1 U990 (.Y(n824), 
	.A(FE_PHN1095_plain_text_94_));
   INVX1 U991 (.Y(n823), 
	.A(FE_PHN2987_plain_text_86_));
   INVX1 U992 (.Y(n822), 
	.A(FE_PHN3000_plain_text_78_));
   INVX1 U993 (.Y(n821), 
	.A(FE_PHN3013_plain_text_70_));
   INVX1 U994 (.Y(n820), 
	.A(FE_PHN2865_plain_text_62_));
   INVX1 U995 (.Y(n819), 
	.A(FE_PHN1196_plain_text_54_));
   INVX1 U996 (.Y(n818), 
	.A(FE_PHN828_plain_text_46_));
   INVX1 U997 (.Y(n817), 
	.A(FE_PHN2022_plain_text_38_));
   INVX1 U998 (.Y(n816), 
	.A(FE_PHN1377_plain_text_30_));
   INVX1 U999 (.Y(n815), 
	.A(FE_PHN3029_plain_text_22_));
   INVX1 U1000 (.Y(n814), 
	.A(FE_PHN3174_plain_text_14_));
   INVX1 U1001 (.Y(n811), 
	.A(FE_PHN1069_plain_text_247_));
   INVX1 U1002 (.Y(n810), 
	.A(FE_PHN1336_plain_text_239_));
   INVX1 U1003 (.Y(n809), 
	.A(FE_PHN1374_plain_text_231_));
   INVX1 U1004 (.Y(n808), 
	.A(FE_PHN3004_plain_text_223_));
   INVX1 U1005 (.Y(n807), 
	.A(FE_PHN1432_plain_text_215_));
   INVX1 U1006 (.Y(n806), 
	.A(FE_PHN1132_plain_text_207_));
   INVX1 U1007 (.Y(n805), 
	.A(FE_PHN2011_plain_text_199_));
   INVX1 U1008 (.Y(n804), 
	.A(FE_PHN3084_plain_text_191_));
   INVX1 U1009 (.Y(n803), 
	.A(FE_PHN1439_plain_text_183_));
   INVX1 U1010 (.Y(n802), 
	.A(FE_PHN3116_plain_text_175_));
   INVX1 U1011 (.Y(n801), 
	.A(FE_PHN1065_plain_text_167_));
   INVX1 U1012 (.Y(n800), 
	.A(FE_PHN3003_plain_text_159_));
   INVX1 U1013 (.Y(n799), 
	.A(FE_PHN2943_plain_text_151_));
   INVX1 U1014 (.Y(n798), 
	.A(FE_PHN2862_plain_text_143_));
   INVX1 U1015 (.Y(n797), 
	.A(FE_PHN2013_plain_text_135_));
   INVX1 U1016 (.Y(n796), 
	.A(FE_PHN1199_plain_text_127_));
   INVX1 U1017 (.Y(n795), 
	.A(FE_PHN2948_plain_text_119_));
   INVX1 U1018 (.Y(n794), 
	.A(FE_PHN1071_plain_text_111_));
   INVX1 U1019 (.Y(n793), 
	.A(FE_PHN1110_plain_text_103_));
   INVX1 U1020 (.Y(n792), 
	.A(FE_PHN1153_plain_text_95_));
   INVX1 U1021 (.Y(n791), 
	.A(FE_PHN1101_plain_text_87_));
   INVX1 U1022 (.Y(n790), 
	.A(FE_PHN3027_plain_text_79_));
   INVX1 U1023 (.Y(n789), 
	.A(FE_PHN1349_plain_text_71_));
   INVX1 U1024 (.Y(n788), 
	.A(FE_PHN1131_plain_text_63_));
   INVX1 U1025 (.Y(n787), 
	.A(FE_PHN1138_plain_text_55_));
   INVX1 U1026 (.Y(n786), 
	.A(FE_PHN1334_plain_text_47_));
   INVX1 U1027 (.Y(n785), 
	.A(FE_PHN2925_plain_text_39_));
   INVX1 U1028 (.Y(n784), 
	.A(FE_PHN1126_plain_text_31_));
   INVX1 U1029 (.Y(n783), 
	.A(FE_PHN1125_plain_text_23_));
   INVX1 U1030 (.Y(n782), 
	.A(FE_PHN2885_plain_text_15_));
   INVX1 U1031 (.Y(n1036), 
	.A(FE_PHN1838_plain_text_248_));
   INVX1 U1032 (.Y(n1004), 
	.A(FE_PHN1218_plain_text_249_));
   INVX1 U1033 (.Y(n972), 
	.A(FE_PHN1242_plain_text_250_));
   INVX1 U1034 (.Y(n940), 
	.A(FE_PHN1250_plain_text_251_));
   INVX1 U1035 (.Y(n908), 
	.A(FE_PHN1240_plain_text_252_));
   INVX1 U1036 (.Y(n876), 
	.A(FE_PHN1228_plain_text_253_));
   INVX1 U1037 (.Y(n844), 
	.A(FE_PHN3087_plain_text_254_));
   INVX1 U1038 (.Y(n812), 
	.A(plain_text[255]));
endmodule

module reg_out (
	clk_48Mhz, 
	reset_n, 
	ready, 
	empty, 
	cipher_text, 
	cipher_byte, 
	cipher_byte_valid, 
	FE_OFN39_reset_n, 
	FE_OFN46_reset_n, 
	FE_OFN50_reset_n, 
	FE_OFN53_reset_n, 
	FE_OFN54_reset_n, 
	FE_OFN55_reset_n, 
	clk_48Mhz__L6_N39, 
	clk_48Mhz__L6_N41, 
	clk_48Mhz__L6_N43, 
	clk_48Mhz__L6_N44, 
	clk_48Mhz__L6_N45, 
	clk_48Mhz__L6_N46, 
	clk_48Mhz__L6_N47);
   input clk_48Mhz;
   input reset_n;
   input ready;
   input empty;
   input [127:0] cipher_text;
   output [7:0] cipher_byte;
   output cipher_byte_valid;
   input FE_OFN39_reset_n;
   input FE_OFN46_reset_n;
   input FE_OFN50_reset_n;
   input FE_OFN53_reset_n;
   input FE_OFN54_reset_n;
   input FE_OFN55_reset_n;
   input clk_48Mhz__L6_N39;
   input clk_48Mhz__L6_N41;
   input clk_48Mhz__L6_N43;
   input clk_48Mhz__L6_N44;
   input clk_48Mhz__L6_N45;
   input clk_48Mhz__L6_N46;
   input clk_48Mhz__L6_N47;

   // Internal wires
   wire FE_PHN5074_n262;
   wire FE_PHN5071_rdy1;
   wire FE_PHN5068_rdy0;
   wire FE_PHN5064_n262;
   wire FE_PHN4962_n368;
   wire FE_PHN4957_n313;
   wire FE_PHN4854_n319;
   wire FE_PHN4666_n320;
   wire FE_PHN4645_n276;
   wire FE_PHN3388_n355;
   wire FE_PHN3378_n363;
   wire FE_PHN3371_cipher_sample_82_;
   wire FE_PHN3365_n283;
   wire FE_PHN3362_n403;
   wire FE_PHN3360_cipher_sample_1_;
   wire FE_PHN3359_n362;
   wire FE_PHN3358_n396;
   wire FE_PHN3356_n196;
   wire FE_PHN3353_cipher_sample_14_;
   wire FE_PHN3351_cipher_sample_93_;
   wire FE_PHN3349_n342;
   wire FE_PHN3345_n424;
   wire FE_PHN3344_n130;
   wire FE_PHN3343_n360;
   wire FE_PHN3342_n303;
   wire FE_PHN3341_n356;
   wire FE_PHN3340_cipher_sample_13_;
   wire FE_PHN3339_n372;
   wire FE_PHN3338_n306;
   wire FE_PHN3335_n371;
   wire FE_PHN3334_n68;
   wire FE_PHN3333_n325;
   wire FE_PHN3332_n334;
   wire FE_PHN3331_n414;
   wire FE_PHN3330_n314;
   wire FE_PHN3329_n407;
   wire FE_PHN3328_n308;
   wire FE_PHN3327_n345;
   wire FE_PHN3326_cipher_sample_30_;
   wire FE_PHN3325_cipher_sample_35_;
   wire FE_PHN3324_n354;
   wire FE_PHN3323_n343;
   wire FE_PHN3322_n340;
   wire FE_PHN3321_n323;
   wire FE_PHN3316_cipher_sample_23_;
   wire FE_PHN3315_n366;
   wire FE_PHN3314_n62;
   wire FE_PHN3313_n358;
   wire FE_PHN3312_cipher_sample_8_;
   wire FE_PHN3310_n286;
   wire FE_PHN3309_cipher_sample_59_;
   wire FE_PHN3308_n330;
   wire FE_PHN3305_n361;
   wire FE_PHN3304_n228;
   wire FE_PHN3302_n353;
   wire FE_PHN3301_cipher_sample_36_;
   wire FE_PHN3296_cipher_sample_52_;
   wire FE_PHN3295_n406;
   wire FE_PHN3294_n337;
   wire FE_PHN3293_n409;
   wire FE_PHN3292_n281;
   wire FE_PHN3290_cipher_sample_41_;
   wire FE_PHN3289_n348;
   wire FE_PHN3288_n311;
   wire FE_PHN3284_n297;
   wire FE_PHN3282_cipher_sample_119_;
   wire FE_PHN3281_cipher_sample_73_;
   wire FE_PHN3278_n316;
   wire FE_PHN3277_cipher_sample_60_;
   wire FE_PHN3276_n329;
   wire FE_PHN3274_n96;
   wire FE_PHN3273_n351;
   wire FE_PHN3272_n294;
   wire FE_PHN3271_n78;
   wire FE_PHN3269_n168;
   wire FE_PHN3268_n290;
   wire FE_PHN3267_n234;
   wire FE_PHN3266_n148;
   wire FE_PHN3265_n194;
   wire FE_PHN3263_n188;
   wire FE_PHN3262_n370;
   wire FE_PHN3261_n418;
   wire FE_PHN3260_n333;
   wire FE_PHN3259_n114;
   wire FE_PHN3256_n74;
   wire FE_PHN3255_n413;
   wire FE_PHN3253_n367;
   wire FE_PHN3252_n301;
   wire FE_PHN3251_n64;
   wire FE_PHN3250_n186;
   wire FE_PHN3249_n305;
   wire FE_PHN3247_n274;
   wire FE_PHN3246_n421;
   wire FE_PHN3245_n309;
   wire FE_PHN3244_cipher_sample_32_;
   wire FE_PHN3243_n357;
   wire FE_PHN3242_n380;
   wire FE_PHN3241_n176;
   wire FE_PHN3240_n289;
   wire FE_PHN3238_cipher_sample_107_;
   wire FE_PHN3237_n282;
   wire FE_PHN3235_n318;
   wire FE_PHN3233_cipher_sample_91_;
   wire FE_PHN3232_n298;
   wire FE_PHN3231_cipher_sample_58_;
   wire FE_PHN3230_n331;
   wire FE_PHN3228_n100;
   wire FE_PHN3227_n335;
   wire FE_PHN3225_n70;
   wire FE_PHN3224_n326;
   wire FE_PHN3223_n76;
   wire FE_PHN3222_n302;
   wire FE_PHN3220_n156;
   wire FE_PHN3219_n369;
   wire FE_PHN3217_cipher_sample_67_;
   wire FE_PHN3216_cipher_sample_102_;
   wire FE_PHN3212_n180;
   wire FE_PHN3211_n273;
   wire FE_PHN3202_n132;
   wire FE_PHN3200_n336;
   wire FE_PHN3193_n312;
   wire FE_PHN3192_n408;
   wire FE_PHN3191_cipher_sample_118_;
   wire FE_PHN3190_n271;
   wire FE_PHN3180_n263;
   wire FE_PHN3179_cipher_sample_122_;
   wire FE_PHN3178_n264;
   wire FE_PHN3177_cipher_sample_123_;
   wire FE_PHN3173_n269;
   wire FE_PHN3161_n268;
   wire FE_PHN3160_n267;
   wire FE_PHN3149_n395;
   wire FE_PHN2993_n376;
   wire FE_PHN2990_n332;
   wire FE_PHN2983_n349;
   wire FE_PHN2982_n327;
   wire FE_PHN2970_n304;
   wire FE_PHN2956_n321;
   wire FE_PHN2955_n315;
   wire FE_PHN2954_n346;
   wire FE_PHN2951_n352;
   wire FE_PHN2947_n373;
   wire FE_PHN2946_n375;
   wire FE_PHN2941_n328;
   wire FE_PHN2936_n322;
   wire FE_PHN2935_n287;
   wire FE_PHN2930_n386;
   wire FE_PHN2927_n284;
   wire FE_PHN2919_cipher_sample_42_;
   wire FE_PHN2918_cipher_sample_2_;
   wire FE_PHN2917_cipher_sample_114_;
   wire FE_PHN2916_cipher_sample_15_;
   wire FE_PHN2915_cipher_sample_12_;
   wire FE_PHN2914_cipher_sample_109_;
   wire FE_PHN2913_n220;
   wire FE_PHN2912_cipher_sample_21_;
   wire FE_PHN2911_n420;
   wire FE_PHN2910_n417;
   wire FE_PHN2909_n106;
   wire FE_PHN2908_n272;
   wire FE_PHN2907_cipher_sample_37_;
   wire FE_PHN2906_cipher_sample_22_;
   wire FE_PHN2905_n350;
   wire FE_PHN2904_n172;
   wire FE_PHN2903_n250;
   wire FE_PHN2902_cipher_sample_94_;
   wire FE_PHN2901_cipher_sample_25_;
   wire FE_PHN2900_n364;
   wire FE_PHN2899_n240;
   wire FE_PHN2898_cipher_sample_0_;
   wire FE_PHN2897_cipher_sample_3_;
   wire FE_PHN2896_cipher_sample_111_;
   wire FE_PHN2895_n138;
   wire FE_PHN2893_cipher_sample_124_;
   wire FE_PHN2892_cipher_sample_127_;
   wire FE_PHN2891_cipher_sample_125_;
   wire FE_PHN2890_cipher_sample_126_;
   wire FE_PHN2849_n293;
   wire FE_PHN2848_n300;
   wire FE_PHN2847_n291;
   wire FE_PHN2846_n389;
   wire FE_PHN2845_n278;
   wire FE_PHN2797_n262;
   wire FE_PHN1458_n263;
   wire FE_PHN1457_n264;
   wire FE_PHN1456_n265;
   wire FE_PHN1455_cipher_sample_120_;
   wire FE_PHN1454_n266;
   wire FE_PHN1449_n269;
   wire FE_PHN1422_n267;
   wire FE_PHN1419_n268;
   wire FE_PHN1380_n392;
   wire FE_PHN1367_n296;
   wire FE_PHN1360_n344;
   wire FE_PHN1353_n342;
   wire FE_PHN1345_n391;
   wire FE_PHN1335_n279;
   wire FE_PHN1299_n307;
   wire FE_PHN1289_n387;
   wire FE_PHN1288_n381;
   wire FE_PHN1284_n365;
   wire FE_PHN1265_n285;
   wire FE_PHN1264_n390;
   wire FE_PHN1262_n292;
   wire FE_PHN1261_n393;
   wire FE_PHN1259_n218;
   wire FE_PHN1258_n120;
   wire FE_PHN1255_n238;
   wire FE_PHN1254_cipher_sample_4_;
   wire FE_PHN1253_n425;
   wire FE_PHN1247_n56;
   wire FE_PHN1237_n144;
   wire FE_PHN1222_n88;
   wire FE_PHN1197_n283;
   wire FE_PHN1172_n396;
   wire FE_PHN1107_n394;
   wire FE_PHN1031_n374;
   wire FE_PHN1030_n376;
   wire FE_PHN1028_n280;
   wire FE_PHN1027_n303;
   wire FE_PHN1026_n366;
   wire FE_PHN1025_n334;
   wire FE_PHN1020_n377;
   wire FE_PHN1019_n351;
   wire FE_PHN1018_n343;
   wire FE_PHN1017_n327;
   wire FE_PHN1013_n368;
   wire FE_PHN1012_n294;
   wire FE_PHN1007_n359;
   wire FE_PHN1004_n272;
   wire FE_PHN1003_n270;
   wire FE_PHN1002_n337;
   wire FE_PHN1001_n375;
   wire FE_PHN987_n310;
   wire FE_PHN985_n328;
   wire FE_PHN978_n281;
   wire FE_PHN967_n369;
   wire FE_PHN952_n295;
   wire FE_PHN951_n273;
   wire FE_PHN946_n302;
   wire FE_PHN941_n335;
   wire FE_PHN931_n326;
   wire FE_PHN927_n367;
   wire FE_PHN926_n288;
   wire FE_PHN925_n336;
   wire FE_PHN920_n278;
   wire FE_PHN918_n271;
   wire FE_PHN887_n355;
   wire FE_PHN885_n275;
   wire FE_PHN881_n363;
   wire FE_PHN879_n356;
   wire FE_PHN878_n324;
   wire FE_PHN877_n347;
   wire FE_PHN876_n372;
   wire FE_PHN873_n319;
   wire FE_PHN872_n345;
   wire FE_PHN871_n338;
   wire FE_PHN869_n306;
   wire FE_PHN868_n341;
   wire FE_PHN867_n353;
   wire FE_PHN866_n360;
   wire FE_PHN865_n325;
   wire FE_PHN863_n388;
   wire FE_PHN862_n332;
   wire FE_PHN859_n339;
   wire FE_PHN858_n379;
   wire FE_PHN857_n397;
   wire FE_PHN856_n340;
   wire FE_PHN855_n333;
   wire FE_PHN854_n330;
   wire FE_PHN853_n320;
   wire FE_PHN852_n276;
   wire FE_PHN851_n384;
   wire FE_PHN850_n297;
   wire FE_PHN849_n286;
   wire FE_PHN848_n316;
   wire FE_PHN847_n370;
   wire FE_PHN846_n301;
   wire FE_PHN845_n299;
   wire FE_PHN844_n358;
   wire FE_PHN843_n371;
   wire FE_PHN842_n385;
   wire FE_PHN841_n290;
   wire FE_PHN840_n277;
   wire FE_PHN839_n298;
   wire FE_PHN838_n361;
   wire FE_PHN836_n318;
   wire FE_PHN834_n382;
   wire FE_PHN833_n331;
   wire FE_PHN832_n311;
   wire FE_PHN831_n305;
   wire FE_PHN826_n312;
   wire FE_PHN825_n383;
   wire FE_PHN818_n349;
   wire FE_PHN816_n362;
   wire FE_PHN815_n314;
   wire FE_PHN814_n313;
   wire FE_PHN813_n323;
   wire FE_PHN809_n317;
   wire FE_PHN805_n348;
   wire FE_PHN804_n354;
   wire FE_PHN801_n289;
   wire FE_PHN799_n321;
   wire FE_PHN795_n346;
   wire FE_PHN793_n329;
   wire FE_PHN790_n308;
   wire FE_PHN787_n380;
   wire FE_PHN784_n322;
   wire FE_PHN781_n357;
   wire FE_PHN778_n378;
   wire FE_PHN761_n386;
   wire FE_PHN759_n284;
   wire FE_PHN729_n304;
   wire FE_PHN725_n352;
   wire FE_PHN697_n373;
   wire FE_PHN695_n274;
   wire FE_PHN693_n364;
   wire FE_PHN690_n287;
   wire FE_PHN687_n309;
   wire FE_PHN685_n350;
   wire FE_PHN636_n315;
   wire FE_PHN634_n300;
   wire FE_PHN630_n389;
   wire FE_PHN629_n291;
   wire FE_PHN505_n395;
   wire FE_PHN445_n282;
   wire FE_PHN358_n293;
   wire FE_PHN124_rdy1;
   wire FE_PHN115_rdy0;
   wire FE_OFN0_n1;
   wire rdy0;
   wire rdy2;
   wire rdy1;
   wire n1;
   wire n5;
   wire n9;
   wire n12;
   wire n15;
   wire n18;
   wire n21;
   wire n24;
   wire n27;
   wire n29;
   wire n31;
   wire n33;
   wire n35;
   wire n37;
   wire n39;
   wire n41;
   wire n43;
   wire n45;
   wire n47;
   wire n49;
   wire n51;
   wire n53;
   wire n55;
   wire n57;
   wire n59;
   wire n61;
   wire n63;
   wire n65;
   wire n67;
   wire n69;
   wire n71;
   wire n73;
   wire n75;
   wire n77;
   wire n79;
   wire n81;
   wire n83;
   wire n85;
   wire n87;
   wire n89;
   wire n91;
   wire n93;
   wire n95;
   wire n97;
   wire n99;
   wire n101;
   wire n103;
   wire n105;
   wire n107;
   wire n109;
   wire n111;
   wire n113;
   wire n115;
   wire n117;
   wire n119;
   wire n121;
   wire n123;
   wire n125;
   wire n127;
   wire n129;
   wire n131;
   wire n133;
   wire n135;
   wire n137;
   wire n139;
   wire n141;
   wire n143;
   wire n145;
   wire n147;
   wire n149;
   wire n151;
   wire n153;
   wire n155;
   wire n157;
   wire n159;
   wire n161;
   wire n163;
   wire n165;
   wire n167;
   wire n169;
   wire n171;
   wire n173;
   wire n175;
   wire n177;
   wire n179;
   wire n181;
   wire n183;
   wire n185;
   wire n187;
   wire n189;
   wire n191;
   wire n193;
   wire n195;
   wire n197;
   wire n199;
   wire n201;
   wire n203;
   wire n205;
   wire n207;
   wire n209;
   wire n211;
   wire n213;
   wire n215;
   wire n217;
   wire n219;
   wire n221;
   wire n223;
   wire n225;
   wire n227;
   wire n229;
   wire n231;
   wire n233;
   wire n235;
   wire n237;
   wire n239;
   wire n241;
   wire n243;
   wire n245;
   wire n247;
   wire n249;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n2;
   wire n4;
   wire n6;
   wire n7;
   wire n8;
   wire n10;
   wire n23;
   wire n25;
   wire n26;
   wire n28;
   wire n30;
   wire n54;
   wire n56;
   wire n58;
   wire n60;
   wire n62;
   wire n64;
   wire n66;
   wire n68;
   wire n70;
   wire n72;
   wire n74;
   wire n76;
   wire n78;
   wire n80;
   wire n82;
   wire n84;
   wire n86;
   wire n88;
   wire n90;
   wire n92;
   wire n94;
   wire n96;
   wire n98;
   wire n100;
   wire n102;
   wire n104;
   wire n106;
   wire n108;
   wire n110;
   wire n112;
   wire n114;
   wire n116;
   wire n118;
   wire n120;
   wire n122;
   wire n124;
   wire n126;
   wire n128;
   wire n130;
   wire n132;
   wire n134;
   wire n136;
   wire n138;
   wire n140;
   wire n142;
   wire n144;
   wire n146;
   wire n148;
   wire n150;
   wire n152;
   wire n154;
   wire n156;
   wire n158;
   wire n160;
   wire n162;
   wire n164;
   wire n166;
   wire n168;
   wire n170;
   wire n172;
   wire n174;
   wire n176;
   wire n178;
   wire n180;
   wire n182;
   wire n184;
   wire n186;
   wire n188;
   wire n190;
   wire n192;
   wire n194;
   wire n196;
   wire n198;
   wire n200;
   wire n202;
   wire n204;
   wire n206;
   wire n208;
   wire n210;
   wire n212;
   wire n214;
   wire n216;
   wire n218;
   wire n220;
   wire n222;
   wire n224;
   wire n226;
   wire n228;
   wire n230;
   wire n232;
   wire n234;
   wire n236;
   wire n238;
   wire n240;
   wire n242;
   wire n244;
   wire n246;
   wire n248;
   wire n250;
   wire n261;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire [127:0] cipher_sample;

   BUFXL FE_PHC5074_n262 (.Y(FE_PHN5074_n262), 
	.A(FE_PHN5064_n262));
   DLY4X1 FE_PHC5071_rdy1 (.Y(FE_PHN5071_rdy1), 
	.A(FE_PHN124_rdy1));
   DLY4X1 FE_PHC5068_rdy0 (.Y(FE_PHN5068_rdy0), 
	.A(FE_PHN115_rdy0));
   CLKBUFX3 FE_PHC5064_n262 (.Y(FE_PHN5064_n262), 
	.A(n262));
   DLY3X1 FE_PHC4962_n368 (.Y(FE_PHN4962_n368), 
	.A(FE_PHN1013_n368));
   DLY4X1 FE_PHC4957_n313 (.Y(FE_PHN4957_n313), 
	.A(n313));
   DLY3X1 FE_PHC4854_n319 (.Y(FE_PHN4854_n319), 
	.A(FE_PHN873_n319));
   DLY4X1 FE_PHC4666_n320 (.Y(FE_PHN4666_n320), 
	.A(FE_PHN853_n320));
   DLY3X1 FE_PHC4645_n276 (.Y(FE_PHN4645_n276), 
	.A(n276));
   DLY3X1 FE_PHC3388_n355 (.Y(FE_PHN3388_n355), 
	.A(FE_PHN887_n355));
   DLY4X1 FE_PHC3378_n363 (.Y(FE_PHN3378_n363), 
	.A(FE_PHN881_n363));
   DLY3X1 FE_PHC3371_cipher_sample_82_ (.Y(FE_PHN3371_cipher_sample_82_), 
	.A(cipher_sample[82]));
   DLY4X1 FE_PHC3365_n283 (.Y(FE_PHN3365_n283), 
	.A(FE_PHN1197_n283));
   DLY3X1 FE_PHC3362_n403 (.Y(FE_PHN3362_n403), 
	.A(n403));
   DLY4X1 FE_PHC3360_cipher_sample_1_ (.Y(FE_PHN3360_cipher_sample_1_), 
	.A(cipher_sample[1]));
   DLY4X1 FE_PHC3359_n362 (.Y(FE_PHN3359_n362), 
	.A(n362));
   DLY4X1 FE_PHC3358_n396 (.Y(FE_PHN3358_n396), 
	.A(n396));
   DLY4X1 FE_PHC3356_n196 (.Y(FE_PHN3356_n196), 
	.A(n196));
   DLY3X1 FE_PHC3353_cipher_sample_14_ (.Y(FE_PHN3353_cipher_sample_14_), 
	.A(cipher_sample[14]));
   DLY3X1 FE_PHC3351_cipher_sample_93_ (.Y(FE_PHN3351_cipher_sample_93_), 
	.A(cipher_sample[93]));
   DLY3X1 FE_PHC3349_n342 (.Y(FE_PHN3349_n342), 
	.A(FE_PHN1353_n342));
   DLY4X1 FE_PHC3345_n424 (.Y(FE_PHN3345_n424), 
	.A(n424));
   DLY4X1 FE_PHC3344_n130 (.Y(FE_PHN3344_n130), 
	.A(n130));
   DLY3X1 FE_PHC3343_n360 (.Y(FE_PHN3343_n360), 
	.A(n360));
   DLY4X1 FE_PHC3342_n303 (.Y(FE_PHN3342_n303), 
	.A(FE_PHN1027_n303));
   DLY4X1 FE_PHC3341_n356 (.Y(FE_PHN3341_n356), 
	.A(FE_PHN879_n356));
   DLY4X1 FE_PHC3340_cipher_sample_13_ (.Y(FE_PHN3340_cipher_sample_13_), 
	.A(cipher_sample[13]));
   DLY4X1 FE_PHC3339_n372 (.Y(FE_PHN3339_n372), 
	.A(n372));
   DLY3X1 FE_PHC3338_n306 (.Y(FE_PHN3338_n306), 
	.A(n306));
   DLY3X1 FE_PHC3335_n371 (.Y(FE_PHN3335_n371), 
	.A(FE_PHN843_n371));
   DLY4X1 FE_PHC3334_n68 (.Y(FE_PHN3334_n68), 
	.A(n68));
   DLY3X1 FE_PHC3333_n325 (.Y(FE_PHN3333_n325), 
	.A(n325));
   DLY3X1 FE_PHC3332_n334 (.Y(FE_PHN3332_n334), 
	.A(FE_PHN1025_n334));
   DLY4X1 FE_PHC3331_n414 (.Y(FE_PHN3331_n414), 
	.A(n414));
   DLY4X1 FE_PHC3330_n314 (.Y(FE_PHN3330_n314), 
	.A(FE_PHN815_n314));
   DLY3X1 FE_PHC3329_n407 (.Y(FE_PHN3329_n407), 
	.A(n407));
   DLY4X1 FE_PHC3328_n308 (.Y(FE_PHN3328_n308), 
	.A(n308));
   DLY4X1 FE_PHC3327_n345 (.Y(FE_PHN3327_n345), 
	.A(FE_PHN872_n345));
   DLY4X1 FE_PHC3326_cipher_sample_30_ (.Y(FE_PHN3326_cipher_sample_30_), 
	.A(cipher_sample[30]));
   DLY4X1 FE_PHC3325_cipher_sample_35_ (.Y(FE_PHN3325_cipher_sample_35_), 
	.A(cipher_sample[35]));
   DLY4X1 FE_PHC3324_n354 (.Y(FE_PHN3324_n354), 
	.A(n354));
   DLY3X1 FE_PHC3323_n343 (.Y(FE_PHN3323_n343), 
	.A(n343));
   DLY3X1 FE_PHC3322_n340 (.Y(FE_PHN3322_n340), 
	.A(FE_PHN856_n340));
   DLY3X1 FE_PHC3321_n323 (.Y(FE_PHN3321_n323), 
	.A(FE_PHN813_n323));
   DLY4X1 FE_PHC3316_cipher_sample_23_ (.Y(FE_PHN3316_cipher_sample_23_), 
	.A(cipher_sample[23]));
   DLY3X1 FE_PHC3315_n366 (.Y(FE_PHN3315_n366), 
	.A(n366));
   DLY4X1 FE_PHC3314_n62 (.Y(FE_PHN3314_n62), 
	.A(n62));
   DLY3X1 FE_PHC3313_n358 (.Y(FE_PHN3313_n358), 
	.A(FE_PHN844_n358));
   DLY4X1 FE_PHC3312_cipher_sample_8_ (.Y(FE_PHN3312_cipher_sample_8_), 
	.A(cipher_sample[8]));
   DLY4X1 FE_PHC3310_n286 (.Y(FE_PHN3310_n286), 
	.A(n286));
   DLY4X1 FE_PHC3309_cipher_sample_59_ (.Y(FE_PHN3309_cipher_sample_59_), 
	.A(cipher_sample[59]));
   DLY3X1 FE_PHC3308_n330 (.Y(FE_PHN3308_n330), 
	.A(FE_PHN854_n330));
   DLY4X1 FE_PHC3305_n361 (.Y(FE_PHN3305_n361), 
	.A(n361));
   DLY3X1 FE_PHC3304_n228 (.Y(FE_PHN3304_n228), 
	.A(n228));
   DLY4X1 FE_PHC3302_n353 (.Y(FE_PHN3302_n353), 
	.A(FE_PHN867_n353));
   DLY4X1 FE_PHC3301_cipher_sample_36_ (.Y(FE_PHN3301_cipher_sample_36_), 
	.A(cipher_sample[36]));
   DLY4X1 FE_PHC3296_cipher_sample_52_ (.Y(FE_PHN3296_cipher_sample_52_), 
	.A(cipher_sample[52]));
   DLY3X1 FE_PHC3295_n406 (.Y(FE_PHN3295_n406), 
	.A(n406));
   DLY3X1 FE_PHC3294_n337 (.Y(FE_PHN3294_n337), 
	.A(n337));
   DLY4X1 FE_PHC3293_n409 (.Y(FE_PHN3293_n409), 
	.A(n409));
   DLY3X1 FE_PHC3292_n281 (.Y(FE_PHN3292_n281), 
	.A(n281));
   DLY4X1 FE_PHC3290_cipher_sample_41_ (.Y(FE_PHN3290_cipher_sample_41_), 
	.A(cipher_sample[41]));
   DLY4X1 FE_PHC3289_n348 (.Y(FE_PHN3289_n348), 
	.A(FE_PHN805_n348));
   DLY4X1 FE_PHC3288_n311 (.Y(FE_PHN3288_n311), 
	.A(n311));
   DLY4X1 FE_PHC3284_n297 (.Y(FE_PHN3284_n297), 
	.A(n297));
   DLY4X1 FE_PHC3282_cipher_sample_119_ (.Y(FE_PHN3282_cipher_sample_119_), 
	.A(cipher_sample[119]));
   DLY4X1 FE_PHC3281_cipher_sample_73_ (.Y(FE_PHN3281_cipher_sample_73_), 
	.A(cipher_sample[73]));
   DLY3X1 FE_PHC3278_n316 (.Y(FE_PHN3278_n316), 
	.A(FE_PHN848_n316));
   DLY4X1 FE_PHC3277_cipher_sample_60_ (.Y(FE_PHN3277_cipher_sample_60_), 
	.A(cipher_sample[60]));
   DLY4X1 FE_PHC3276_n329 (.Y(FE_PHN3276_n329), 
	.A(n329));
   DLY4X1 FE_PHC3274_n96 (.Y(FE_PHN3274_n96), 
	.A(n96));
   DLY4X1 FE_PHC3273_n351 (.Y(FE_PHN3273_n351), 
	.A(FE_PHN1019_n351));
   DLY4X1 FE_PHC3272_n294 (.Y(FE_PHN3272_n294), 
	.A(FE_PHN1012_n294));
   DLY4X1 FE_PHC3271_n78 (.Y(FE_PHN3271_n78), 
	.A(n78));
   DLY4X1 FE_PHC3269_n168 (.Y(FE_PHN3269_n168), 
	.A(n168));
   DLY4X1 FE_PHC3268_n290 (.Y(FE_PHN3268_n290), 
	.A(n290));
   DLY4X1 FE_PHC3267_n234 (.Y(FE_PHN3267_n234), 
	.A(n234));
   DLY4X1 FE_PHC3266_n148 (.Y(FE_PHN3266_n148), 
	.A(n148));
   DLY4X1 FE_PHC3265_n194 (.Y(FE_PHN3265_n194), 
	.A(n194));
   DLY4X1 FE_PHC3263_n188 (.Y(FE_PHN3263_n188), 
	.A(n188));
   DLY4X1 FE_PHC3262_n370 (.Y(FE_PHN3262_n370), 
	.A(n370));
   DLY4X1 FE_PHC3261_n418 (.Y(FE_PHN3261_n418), 
	.A(n418));
   DLY4X1 FE_PHC3260_n333 (.Y(FE_PHN3260_n333), 
	.A(FE_PHN855_n333));
   DLY4X1 FE_PHC3259_n114 (.Y(FE_PHN3259_n114), 
	.A(n114));
   DLY4X1 FE_PHC3256_n74 (.Y(FE_PHN3256_n74), 
	.A(n74));
   DLY4X1 FE_PHC3255_n413 (.Y(FE_PHN3255_n413), 
	.A(n413));
   DLY4X1 FE_PHC3253_n367 (.Y(FE_PHN3253_n367), 
	.A(n367));
   DLY4X1 FE_PHC3252_n301 (.Y(FE_PHN3252_n301), 
	.A(FE_PHN846_n301));
   DLY3X1 FE_PHC3251_n64 (.Y(FE_PHN3251_n64), 
	.A(n64));
   DLY4X1 FE_PHC3250_n186 (.Y(FE_PHN3250_n186), 
	.A(n186));
   DLY4X1 FE_PHC3249_n305 (.Y(FE_PHN3249_n305), 
	.A(n305));
   DLY4X1 FE_PHC3247_n274 (.Y(FE_PHN3247_n274), 
	.A(n274));
   DLY4X1 FE_PHC3246_n421 (.Y(FE_PHN3246_n421), 
	.A(n421));
   DLY4X1 FE_PHC3245_n309 (.Y(FE_PHN3245_n309), 
	.A(n309));
   DLY4X1 FE_PHC3244_cipher_sample_32_ (.Y(FE_PHN3244_cipher_sample_32_), 
	.A(cipher_sample[32]));
   DLY4X1 FE_PHC3243_n357 (.Y(FE_PHN3243_n357), 
	.A(n357));
   DLY4X1 FE_PHC3242_n380 (.Y(FE_PHN3242_n380), 
	.A(n380));
   DLY4X1 FE_PHC3241_n176 (.Y(FE_PHN3241_n176), 
	.A(n176));
   DLY4X1 FE_PHC3240_n289 (.Y(FE_PHN3240_n289), 
	.A(n289));
   DLY4X1 FE_PHC3238_cipher_sample_107_ (.Y(FE_PHN3238_cipher_sample_107_), 
	.A(cipher_sample[107]));
   DLY4X1 FE_PHC3237_n282 (.Y(FE_PHN3237_n282), 
	.A(n282));
   DLY4X1 FE_PHC3235_n318 (.Y(FE_PHN3235_n318), 
	.A(n318));
   DLY4X1 FE_PHC3233_cipher_sample_91_ (.Y(FE_PHN3233_cipher_sample_91_), 
	.A(cipher_sample[91]));
   DLY4X1 FE_PHC3232_n298 (.Y(FE_PHN3232_n298), 
	.A(n298));
   DLY4X1 FE_PHC3231_cipher_sample_58_ (.Y(FE_PHN3231_cipher_sample_58_), 
	.A(cipher_sample[58]));
   DLY4X1 FE_PHC3230_n331 (.Y(FE_PHN3230_n331), 
	.A(n331));
   DLY4X1 FE_PHC3228_n100 (.Y(FE_PHN3228_n100), 
	.A(n100));
   DLY4X1 FE_PHC3227_n335 (.Y(FE_PHN3227_n335), 
	.A(n335));
   DLY4X1 FE_PHC3225_n70 (.Y(FE_PHN3225_n70), 
	.A(n70));
   DLY4X1 FE_PHC3224_n326 (.Y(FE_PHN3224_n326), 
	.A(n326));
   DLY4X1 FE_PHC3223_n76 (.Y(FE_PHN3223_n76), 
	.A(n76));
   DLY4X1 FE_PHC3222_n302 (.Y(FE_PHN3222_n302), 
	.A(n302));
   DLY4X1 FE_PHC3220_n156 (.Y(FE_PHN3220_n156), 
	.A(n156));
   DLY4X1 FE_PHC3219_n369 (.Y(FE_PHN3219_n369), 
	.A(n369));
   DLY4X1 FE_PHC3217_cipher_sample_67_ (.Y(FE_PHN3217_cipher_sample_67_), 
	.A(cipher_sample[67]));
   DLY4X1 FE_PHC3216_cipher_sample_102_ (.Y(FE_PHN3216_cipher_sample_102_), 
	.A(cipher_sample[102]));
   DLY4X1 FE_PHC3212_n180 (.Y(FE_PHN3212_n180), 
	.A(n180));
   DLY4X1 FE_PHC3211_n273 (.Y(FE_PHN3211_n273), 
	.A(n273));
   DLY4X1 FE_PHC3202_n132 (.Y(FE_PHN3202_n132), 
	.A(n132));
   DLY4X1 FE_PHC3200_n336 (.Y(FE_PHN3200_n336), 
	.A(n336));
   DLY4X1 FE_PHC3193_n312 (.Y(FE_PHN3193_n312), 
	.A(n312));
   DLY4X1 FE_PHC3192_n408 (.Y(FE_PHN3192_n408), 
	.A(n408));
   DLY4X1 FE_PHC3191_cipher_sample_118_ (.Y(FE_PHN3191_cipher_sample_118_), 
	.A(cipher_sample[118]));
   DLY4X1 FE_PHC3190_n271 (.Y(FE_PHN3190_n271), 
	.A(n271));
   DLY2X1 FE_PHC3180_n263 (.Y(FE_PHN3180_n263), 
	.A(n263));
   DLY2X1 FE_PHC3179_cipher_sample_122_ (.Y(FE_PHN3179_cipher_sample_122_), 
	.A(cipher_sample[122]));
   DLY2X1 FE_PHC3178_n264 (.Y(FE_PHN3178_n264), 
	.A(n264));
   DLY2X1 FE_PHC3177_cipher_sample_123_ (.Y(FE_PHN3177_cipher_sample_123_), 
	.A(cipher_sample[123]));
   DLY4X1 FE_PHC3173_n269 (.Y(FE_PHN3173_n269), 
	.A(n269));
   DLY4X1 FE_PHC3161_n268 (.Y(FE_PHN3161_n268), 
	.A(n268));
   DLY4X1 FE_PHC3160_n267 (.Y(FE_PHN3160_n267), 
	.A(n267));
   DLY3X1 FE_PHC3149_n395 (.Y(FE_PHN3149_n395), 
	.A(n395));
   DLY4X1 FE_PHC2993_n376 (.Y(FE_PHN2993_n376), 
	.A(n376));
   DLY4X1 FE_PHC2990_n332 (.Y(FE_PHN2990_n332), 
	.A(FE_PHN862_n332));
   DLY4X1 FE_PHC2983_n349 (.Y(FE_PHN2983_n349), 
	.A(n349));
   DLY3X1 FE_PHC2982_n327 (.Y(FE_PHN2982_n327), 
	.A(n327));
   DLY4X1 FE_PHC2970_n304 (.Y(FE_PHN2970_n304), 
	.A(n304));
   DLY4X1 FE_PHC2956_n321 (.Y(FE_PHN2956_n321), 
	.A(n321));
   DLY4X1 FE_PHC2955_n315 (.Y(FE_PHN2955_n315), 
	.A(n315));
   DLY4X1 FE_PHC2954_n346 (.Y(FE_PHN2954_n346), 
	.A(n346));
   DLY3X1 FE_PHC2951_n352 (.Y(FE_PHN2951_n352), 
	.A(n352));
   DLY4X1 FE_PHC2947_n373 (.Y(FE_PHN2947_n373), 
	.A(n373));
   DLY4X1 FE_PHC2946_n375 (.Y(FE_PHN2946_n375), 
	.A(n375));
   DLY4X1 FE_PHC2941_n328 (.Y(FE_PHN2941_n328), 
	.A(n328));
   DLY4X1 FE_PHC2936_n322 (.Y(FE_PHN2936_n322), 
	.A(n322));
   DLY4X1 FE_PHC2935_n287 (.Y(FE_PHN2935_n287), 
	.A(n287));
   DLY4X1 FE_PHC2930_n386 (.Y(FE_PHN2930_n386), 
	.A(n386));
   DLY4X1 FE_PHC2927_n284 (.Y(FE_PHN2927_n284), 
	.A(n284));
   DLY4X1 FE_PHC2919_cipher_sample_42_ (.Y(FE_PHN2919_cipher_sample_42_), 
	.A(cipher_sample[42]));
   DLY4X1 FE_PHC2918_cipher_sample_2_ (.Y(FE_PHN2918_cipher_sample_2_), 
	.A(cipher_sample[2]));
   DLY4X1 FE_PHC2917_cipher_sample_114_ (.Y(FE_PHN2917_cipher_sample_114_), 
	.A(cipher_sample[114]));
   DLY4X1 FE_PHC2916_cipher_sample_15_ (.Y(FE_PHN2916_cipher_sample_15_), 
	.A(cipher_sample[15]));
   DLY4X1 FE_PHC2915_cipher_sample_12_ (.Y(FE_PHN2915_cipher_sample_12_), 
	.A(cipher_sample[12]));
   DLY4X1 FE_PHC2914_cipher_sample_109_ (.Y(FE_PHN2914_cipher_sample_109_), 
	.A(cipher_sample[109]));
   DLY3X1 FE_PHC2913_n220 (.Y(FE_PHN2913_n220), 
	.A(n220));
   DLY4X1 FE_PHC2912_cipher_sample_21_ (.Y(FE_PHN2912_cipher_sample_21_), 
	.A(cipher_sample[21]));
   DLY3X1 FE_PHC2911_n420 (.Y(FE_PHN2911_n420), 
	.A(n420));
   DLY4X1 FE_PHC2910_n417 (.Y(FE_PHN2910_n417), 
	.A(n417));
   DLY4X1 FE_PHC2909_n106 (.Y(FE_PHN2909_n106), 
	.A(n106));
   DLY4X1 FE_PHC2908_n272 (.Y(FE_PHN2908_n272), 
	.A(FE_PHN1004_n272));
   DLY4X1 FE_PHC2907_cipher_sample_37_ (.Y(FE_PHN2907_cipher_sample_37_), 
	.A(cipher_sample[37]));
   DLY4X1 FE_PHC2906_cipher_sample_22_ (.Y(FE_PHN2906_cipher_sample_22_), 
	.A(cipher_sample[22]));
   DLY4X1 FE_PHC2905_n350 (.Y(FE_PHN2905_n350), 
	.A(n350));
   DLY4X1 FE_PHC2904_n172 (.Y(FE_PHN2904_n172), 
	.A(n172));
   DLY4X1 FE_PHC2903_n250 (.Y(FE_PHN2903_n250), 
	.A(n250));
   DLY4X1 FE_PHC2902_cipher_sample_94_ (.Y(FE_PHN2902_cipher_sample_94_), 
	.A(cipher_sample[94]));
   DLY4X1 FE_PHC2901_cipher_sample_25_ (.Y(FE_PHN2901_cipher_sample_25_), 
	.A(cipher_sample[25]));
   DLY4X1 FE_PHC2900_n364 (.Y(FE_PHN2900_n364), 
	.A(n364));
   DLY4X1 FE_PHC2899_n240 (.Y(FE_PHN2899_n240), 
	.A(n240));
   DLY4X1 FE_PHC2898_cipher_sample_0_ (.Y(FE_PHN2898_cipher_sample_0_), 
	.A(cipher_sample[0]));
   DLY4X1 FE_PHC2897_cipher_sample_3_ (.Y(FE_PHN2897_cipher_sample_3_), 
	.A(cipher_sample[3]));
   DLY4X1 FE_PHC2896_cipher_sample_111_ (.Y(FE_PHN2896_cipher_sample_111_), 
	.A(cipher_sample[111]));
   DLY4X1 FE_PHC2895_n138 (.Y(FE_PHN2895_n138), 
	.A(n138));
   DLY3X1 FE_PHC2893_cipher_sample_124_ (.Y(FE_PHN2893_cipher_sample_124_), 
	.A(cipher_sample[124]));
   DLY4X1 FE_PHC2892_cipher_sample_127_ (.Y(FE_PHN2892_cipher_sample_127_), 
	.A(cipher_sample[127]));
   DLY4X1 FE_PHC2891_cipher_sample_125_ (.Y(FE_PHN2891_cipher_sample_125_), 
	.A(cipher_sample[125]));
   DLY4X1 FE_PHC2890_cipher_sample_126_ (.Y(FE_PHN2890_cipher_sample_126_), 
	.A(cipher_sample[126]));
   DLY4X1 FE_PHC2849_n293 (.Y(FE_PHN2849_n293), 
	.A(n293));
   DLY3X1 FE_PHC2848_n300 (.Y(FE_PHN2848_n300), 
	.A(n300));
   DLY4X1 FE_PHC2847_n291 (.Y(FE_PHN2847_n291), 
	.A(n291));
   DLY4X1 FE_PHC2846_n389 (.Y(FE_PHN2846_n389), 
	.A(n389));
   DLY4X1 FE_PHC2845_n278 (.Y(FE_PHN2845_n278), 
	.A(n278));
   DLY4X1 FE_PHC2797_n262 (.Y(FE_PHN2797_n262), 
	.A(FE_PHN5074_n262));
   DLY4X1 FE_PHC1458_n263 (.Y(FE_PHN1458_n263), 
	.A(FE_PHN3180_n263));
   DLY4X1 FE_PHC1457_n264 (.Y(FE_PHN1457_n264), 
	.A(FE_PHN3178_n264));
   DLY4X1 FE_PHC1456_n265 (.Y(FE_PHN1456_n265), 
	.A(n265));
   DLY4X1 FE_PHC1455_cipher_sample_120_ (.Y(FE_PHN1455_cipher_sample_120_), 
	.A(cipher_sample[120]));
   DLY4X1 FE_PHC1454_n266 (.Y(FE_PHN1454_n266), 
	.A(n266));
   DLY4X1 FE_PHC1449_n269 (.Y(FE_PHN1449_n269), 
	.A(FE_PHN3173_n269));
   DLY4X1 FE_PHC1422_n267 (.Y(FE_PHN1422_n267), 
	.A(FE_PHN3160_n267));
   DLY4X1 FE_PHC1419_n268 (.Y(FE_PHN1419_n268), 
	.A(FE_PHN3161_n268));
   DLY4X1 FE_PHC1380_n392 (.Y(FE_PHN1380_n392), 
	.A(n392));
   DLY4X1 FE_PHC1367_n296 (.Y(FE_PHN1367_n296), 
	.A(n296));
   DLY4X1 FE_PHC1360_n344 (.Y(FE_PHN1360_n344), 
	.A(n344));
   DLY4X1 FE_PHC1353_n342 (.Y(FE_PHN1353_n342), 
	.A(n342));
   DLY4X1 FE_PHC1345_n391 (.Y(FE_PHN1345_n391), 
	.A(n391));
   DLY4X1 FE_PHC1335_n279 (.Y(FE_PHN1335_n279), 
	.A(n279));
   DLY4X1 FE_PHC1299_n307 (.Y(FE_PHN1299_n307), 
	.A(n307));
   DLY4X1 FE_PHC1289_n387 (.Y(FE_PHN1289_n387), 
	.A(n387));
   DLY4X1 FE_PHC1288_n381 (.Y(FE_PHN1288_n381), 
	.A(n381));
   DLY4X1 FE_PHC1284_n365 (.Y(FE_PHN1284_n365), 
	.A(n365));
   DLY4X1 FE_PHC1265_n285 (.Y(FE_PHN1265_n285), 
	.A(n285));
   DLY4X1 FE_PHC1264_n390 (.Y(FE_PHN1264_n390), 
	.A(n390));
   DLY4X1 FE_PHC1262_n292 (.Y(FE_PHN1262_n292), 
	.A(n292));
   DLY4X1 FE_PHC1261_n393 (.Y(FE_PHN1261_n393), 
	.A(n393));
   DLY4X1 FE_PHC1259_n218 (.Y(FE_PHN1259_n218), 
	.A(n218));
   DLY4X1 FE_PHC1258_n120 (.Y(FE_PHN1258_n120), 
	.A(n120));
   DLY4X1 FE_PHC1255_n238 (.Y(FE_PHN1255_n238), 
	.A(n238));
   DLY4X1 FE_PHC1254_cipher_sample_4_ (.Y(FE_PHN1254_cipher_sample_4_), 
	.A(cipher_sample[4]));
   DLY4X1 FE_PHC1253_n425 (.Y(FE_PHN1253_n425), 
	.A(n425));
   DLY4X1 FE_PHC1247_n56 (.Y(FE_PHN1247_n56), 
	.A(n56));
   DLY4X1 FE_PHC1237_n144 (.Y(FE_PHN1237_n144), 
	.A(n144));
   DLY4X1 FE_PHC1222_n88 (.Y(FE_PHN1222_n88), 
	.A(n88));
   DLY4X1 FE_PHC1197_n283 (.Y(FE_PHN1197_n283), 
	.A(n283));
   DLY4X1 FE_PHC1172_n396 (.Y(FE_PHN1172_n396), 
	.A(FE_PHN3358_n396));
   DLY4X1 FE_PHC1107_n394 (.Y(FE_PHN1107_n394), 
	.A(n394));
   DLY4X1 FE_PHC1031_n374 (.Y(FE_PHN1031_n374), 
	.A(n374));
   DLY4X1 FE_PHC1030_n376 (.Y(FE_PHN1030_n376), 
	.A(FE_PHN2993_n376));
   DLY4X1 FE_PHC1028_n280 (.Y(FE_PHN1028_n280), 
	.A(n280));
   DLY4X1 FE_PHC1027_n303 (.Y(FE_PHN1027_n303), 
	.A(n303));
   DLY4X1 FE_PHC1026_n366 (.Y(FE_PHN1026_n366), 
	.A(FE_PHN3315_n366));
   DLY4X1 FE_PHC1025_n334 (.Y(FE_PHN1025_n334), 
	.A(n334));
   DLY4X1 FE_PHC1020_n377 (.Y(FE_PHN1020_n377), 
	.A(n377));
   DLY4X1 FE_PHC1019_n351 (.Y(FE_PHN1019_n351), 
	.A(n351));
   DLY4X1 FE_PHC1018_n343 (.Y(FE_PHN1018_n343), 
	.A(FE_PHN3323_n343));
   DLY4X1 FE_PHC1017_n327 (.Y(FE_PHN1017_n327), 
	.A(FE_PHN2982_n327));
   DLY4X1 FE_PHC1013_n368 (.Y(FE_PHN1013_n368), 
	.A(n368));
   DLY4X1 FE_PHC1012_n294 (.Y(FE_PHN1012_n294), 
	.A(n294));
   DLY4X1 FE_PHC1007_n359 (.Y(FE_PHN1007_n359), 
	.A(n359));
   DLY4X1 FE_PHC1004_n272 (.Y(FE_PHN1004_n272), 
	.A(n272));
   DLY4X1 FE_PHC1003_n270 (.Y(FE_PHN1003_n270), 
	.A(n270));
   DLY4X1 FE_PHC1002_n337 (.Y(FE_PHN1002_n337), 
	.A(FE_PHN3294_n337));
   DLY4X1 FE_PHC1001_n375 (.Y(FE_PHN1001_n375), 
	.A(FE_PHN2946_n375));
   DLY4X1 FE_PHC987_n310 (.Y(FE_PHN987_n310), 
	.A(n310));
   DLY4X1 FE_PHC985_n328 (.Y(FE_PHN985_n328), 
	.A(FE_PHN2941_n328));
   DLY4X1 FE_PHC978_n281 (.Y(FE_PHN978_n281), 
	.A(FE_PHN3292_n281));
   DLY4X1 FE_PHC967_n369 (.Y(FE_PHN967_n369), 
	.A(FE_PHN3219_n369));
   DLY4X1 FE_PHC952_n295 (.Y(FE_PHN952_n295), 
	.A(n295));
   DLY4X1 FE_PHC951_n273 (.Y(FE_PHN951_n273), 
	.A(FE_PHN3211_n273));
   DLY4X1 FE_PHC946_n302 (.Y(FE_PHN946_n302), 
	.A(FE_PHN3222_n302));
   DLY4X1 FE_PHC941_n335 (.Y(FE_PHN941_n335), 
	.A(FE_PHN3227_n335));
   DLY4X1 FE_PHC931_n326 (.Y(FE_PHN931_n326), 
	.A(FE_PHN3224_n326));
   DLY4X1 FE_PHC927_n367 (.Y(FE_PHN927_n367), 
	.A(FE_PHN3253_n367));
   DLY4X1 FE_PHC926_n288 (.Y(FE_PHN926_n288), 
	.A(n288));
   DLY4X1 FE_PHC925_n336 (.Y(FE_PHN925_n336), 
	.A(FE_PHN3200_n336));
   DLY4X1 FE_PHC920_n278 (.Y(FE_PHN920_n278), 
	.A(FE_PHN2845_n278));
   DLY4X1 FE_PHC918_n271 (.Y(FE_PHN918_n271), 
	.A(FE_PHN3190_n271));
   DLY4X1 FE_PHC887_n355 (.Y(FE_PHN887_n355), 
	.A(n355));
   DLY4X1 FE_PHC885_n275 (.Y(FE_PHN885_n275), 
	.A(n275));
   DLY4X1 FE_PHC881_n363 (.Y(FE_PHN881_n363), 
	.A(n363));
   DLY4X1 FE_PHC879_n356 (.Y(FE_PHN879_n356), 
	.A(n356));
   DLY4X1 FE_PHC878_n324 (.Y(FE_PHN878_n324), 
	.A(n324));
   DLY4X1 FE_PHC877_n347 (.Y(FE_PHN877_n347), 
	.A(n347));
   DLY4X1 FE_PHC876_n372 (.Y(FE_PHN876_n372), 
	.A(FE_PHN3339_n372));
   DLY4X1 FE_PHC873_n319 (.Y(FE_PHN873_n319), 
	.A(n319));
   DLY4X1 FE_PHC872_n345 (.Y(FE_PHN872_n345), 
	.A(n345));
   DLY4X1 FE_PHC871_n338 (.Y(FE_PHN871_n338), 
	.A(n338));
   DLY4X1 FE_PHC869_n306 (.Y(FE_PHN869_n306), 
	.A(FE_PHN3338_n306));
   DLY4X1 FE_PHC868_n341 (.Y(FE_PHN868_n341), 
	.A(n341));
   DLY4X1 FE_PHC867_n353 (.Y(FE_PHN867_n353), 
	.A(n353));
   DLY4X1 FE_PHC866_n360 (.Y(FE_PHN866_n360), 
	.A(FE_PHN3343_n360));
   DLY4X1 FE_PHC865_n325 (.Y(FE_PHN865_n325), 
	.A(FE_PHN3333_n325));
   DLY4X1 FE_PHC863_n388 (.Y(FE_PHN863_n388), 
	.A(n388));
   DLY4X1 FE_PHC862_n332 (.Y(FE_PHN862_n332), 
	.A(n332));
   DLY4X1 FE_PHC859_n339 (.Y(FE_PHN859_n339), 
	.A(n339));
   DLY4X1 FE_PHC858_n379 (.Y(FE_PHN858_n379), 
	.A(n379));
   DLY4X1 FE_PHC857_n397 (.Y(FE_PHN857_n397), 
	.A(n397));
   DLY4X1 FE_PHC856_n340 (.Y(FE_PHN856_n340), 
	.A(n340));
   DLY4X1 FE_PHC855_n333 (.Y(FE_PHN855_n333), 
	.A(n333));
   DLY4X1 FE_PHC854_n330 (.Y(FE_PHN854_n330), 
	.A(n330));
   DLY4X1 FE_PHC853_n320 (.Y(FE_PHN853_n320), 
	.A(n320));
   DLY4X1 FE_PHC852_n276 (.Y(FE_PHN852_n276), 
	.A(FE_PHN4645_n276));
   DLY4X1 FE_PHC851_n384 (.Y(FE_PHN851_n384), 
	.A(n384));
   DLY4X1 FE_PHC850_n297 (.Y(FE_PHN850_n297), 
	.A(FE_PHN3284_n297));
   DLY4X1 FE_PHC849_n286 (.Y(FE_PHN849_n286), 
	.A(FE_PHN3310_n286));
   DLY4X1 FE_PHC848_n316 (.Y(FE_PHN848_n316), 
	.A(n316));
   DLY4X1 FE_PHC847_n370 (.Y(FE_PHN847_n370), 
	.A(FE_PHN3262_n370));
   DLY4X1 FE_PHC846_n301 (.Y(FE_PHN846_n301), 
	.A(n301));
   DLY4X1 FE_PHC845_n299 (.Y(FE_PHN845_n299), 
	.A(n299));
   DLY4X1 FE_PHC844_n358 (.Y(FE_PHN844_n358), 
	.A(n358));
   DLY4X1 FE_PHC843_n371 (.Y(FE_PHN843_n371), 
	.A(n371));
   DLY4X1 FE_PHC842_n385 (.Y(FE_PHN842_n385), 
	.A(n385));
   DLY4X1 FE_PHC841_n290 (.Y(FE_PHN841_n290), 
	.A(FE_PHN3268_n290));
   DLY4X1 FE_PHC840_n277 (.Y(FE_PHN840_n277), 
	.A(n277));
   DLY4X1 FE_PHC839_n298 (.Y(FE_PHN839_n298), 
	.A(FE_PHN3232_n298));
   DLY4X1 FE_PHC838_n361 (.Y(FE_PHN838_n361), 
	.A(FE_PHN3305_n361));
   DLY4X1 FE_PHC836_n318 (.Y(FE_PHN836_n318), 
	.A(FE_PHN3235_n318));
   DLY4X1 FE_PHC834_n382 (.Y(FE_PHN834_n382), 
	.A(n382));
   DLY4X1 FE_PHC833_n331 (.Y(FE_PHN833_n331), 
	.A(FE_PHN3230_n331));
   DLY4X1 FE_PHC832_n311 (.Y(FE_PHN832_n311), 
	.A(FE_PHN3288_n311));
   DLY4X1 FE_PHC831_n305 (.Y(FE_PHN831_n305), 
	.A(FE_PHN3249_n305));
   DLY4X1 FE_PHC826_n312 (.Y(FE_PHN826_n312), 
	.A(FE_PHN3193_n312));
   DLY4X1 FE_PHC825_n383 (.Y(FE_PHN825_n383), 
	.A(n383));
   DLY4X1 FE_PHC818_n349 (.Y(FE_PHN818_n349), 
	.A(FE_PHN2983_n349));
   DLY4X1 FE_PHC816_n362 (.Y(FE_PHN816_n362), 
	.A(FE_PHN3359_n362));
   DLY4X1 FE_PHC815_n314 (.Y(FE_PHN815_n314), 
	.A(n314));
   DLY4X1 FE_PHC814_n313 (.Y(FE_PHN814_n313), 
	.A(FE_PHN4957_n313));
   DLY4X1 FE_PHC813_n323 (.Y(FE_PHN813_n323), 
	.A(n323));
   DLY4X1 FE_PHC809_n317 (.Y(FE_PHN809_n317), 
	.A(n317));
   DLY4X1 FE_PHC805_n348 (.Y(FE_PHN805_n348), 
	.A(n348));
   DLY4X1 FE_PHC804_n354 (.Y(FE_PHN804_n354), 
	.A(FE_PHN3324_n354));
   DLY4X1 FE_PHC801_n289 (.Y(FE_PHN801_n289), 
	.A(FE_PHN3240_n289));
   DLY4X1 FE_PHC799_n321 (.Y(FE_PHN799_n321), 
	.A(FE_PHN2956_n321));
   DLY4X1 FE_PHC795_n346 (.Y(FE_PHN795_n346), 
	.A(FE_PHN2954_n346));
   DLY4X1 FE_PHC793_n329 (.Y(FE_PHN793_n329), 
	.A(FE_PHN3276_n329));
   DLY4X1 FE_PHC790_n308 (.Y(FE_PHN790_n308), 
	.A(FE_PHN3328_n308));
   DLY4X1 FE_PHC787_n380 (.Y(FE_PHN787_n380), 
	.A(FE_PHN3242_n380));
   DLY4X1 FE_PHC784_n322 (.Y(FE_PHN784_n322), 
	.A(FE_PHN2936_n322));
   DLY4X1 FE_PHC781_n357 (.Y(FE_PHN781_n357), 
	.A(FE_PHN3243_n357));
   DLY4X1 FE_PHC778_n378 (.Y(FE_PHN778_n378), 
	.A(n378));
   DLY4X1 FE_PHC761_n386 (.Y(FE_PHN761_n386), 
	.A(FE_PHN2930_n386));
   DLY4X1 FE_PHC759_n284 (.Y(FE_PHN759_n284), 
	.A(FE_PHN2927_n284));
   DLY4X1 FE_PHC729_n304 (.Y(FE_PHN729_n304), 
	.A(FE_PHN2970_n304));
   DLY4X1 FE_PHC725_n352 (.Y(FE_PHN725_n352), 
	.A(FE_PHN2951_n352));
   DLY4X1 FE_PHC697_n373 (.Y(FE_PHN697_n373), 
	.A(FE_PHN2947_n373));
   DLY4X1 FE_PHC695_n274 (.Y(FE_PHN695_n274), 
	.A(FE_PHN3247_n274));
   DLY4X1 FE_PHC693_n364 (.Y(FE_PHN693_n364), 
	.A(FE_PHN2900_n364));
   DLY4X1 FE_PHC690_n287 (.Y(FE_PHN690_n287), 
	.A(FE_PHN2935_n287));
   DLY4X1 FE_PHC687_n309 (.Y(FE_PHN687_n309), 
	.A(FE_PHN3245_n309));
   DLY4X1 FE_PHC685_n350 (.Y(FE_PHN685_n350), 
	.A(FE_PHN2905_n350));
   DLY4X1 FE_PHC636_n315 (.Y(FE_PHN636_n315), 
	.A(FE_PHN2955_n315));
   DLY4X1 FE_PHC634_n300 (.Y(FE_PHN634_n300), 
	.A(FE_PHN2848_n300));
   DLY4X1 FE_PHC630_n389 (.Y(FE_PHN630_n389), 
	.A(FE_PHN2846_n389));
   DLY4X1 FE_PHC629_n291 (.Y(FE_PHN629_n291), 
	.A(FE_PHN2847_n291));
   DLY4X1 FE_PHC505_n395 (.Y(FE_PHN505_n395), 
	.A(FE_PHN3149_n395));
   DLY4X1 FE_PHC445_n282 (.Y(FE_PHN445_n282), 
	.A(FE_PHN3237_n282));
   DLY4X1 FE_PHC358_n293 (.Y(FE_PHN358_n293), 
	.A(FE_PHN2849_n293));
   DLY4X1 FE_PHC124_rdy1 (.Y(FE_PHN124_rdy1), 
	.A(rdy1));
   DLY4X1 FE_PHC115_rdy0 (.Y(FE_PHN115_rdy0), 
	.A(rdy0));
   CLKBUFX2 FE_OFC0_n1 (.Y(FE_OFN0_n1), 
	.A(n1));
   DFFRHQX1 cipher_sample_reg_7_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[7]), 
	.D(FE_PHN1264_n390), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_15_ (.RN(reset_n), 
	.Q(cipher_sample[15]), 
	.D(FE_PHN834_n382), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_23_ (.RN(reset_n), 
	.Q(cipher_sample[23]), 
	.D(FE_PHN1031_n374), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_31_ (.RN(reset_n), 
	.Q(cipher_sample[31]), 
	.D(FE_PHN1026_n366), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_39_ (.RN(reset_n), 
	.Q(cipher_sample[39]), 
	.D(FE_PHN3313_n358), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_47_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[47]), 
	.D(FE_PHN685_n350), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_55_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[55]), 
	.D(FE_PHN3349_n342), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_63_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[63]), 
	.D(FE_PHN3332_n334), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_71_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[71]), 
	.D(FE_PHN931_n326), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_79_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[79]), 
	.D(FE_PHN836_n318), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_87_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[87]), 
	.D(FE_PHN987_n310), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_95_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[95]), 
	.D(FE_PHN946_n302), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_103_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[103]), 
	.D(FE_PHN3272_n294), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_111_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[111]), 
	.D(FE_PHN849_n286), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_119_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[119]), 
	.D(FE_PHN920_n278), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_127_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[127]), 
	.D(FE_PHN1003_n270), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_6_ (.RN(reset_n), 
	.Q(cipher_sample[6]), 
	.D(FE_PHN1345_n391), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_14_ (.RN(reset_n), 
	.Q(cipher_sample[14]), 
	.D(FE_PHN825_n383), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_22_ (.RN(reset_n), 
	.Q(cipher_sample[22]), 
	.D(FE_PHN1001_n375), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 cipher_sample_reg_30_ (.RN(reset_n), 
	.Q(cipher_sample[30]), 
	.D(FE_PHN927_n367), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 cipher_sample_reg_38_ (.RN(reset_n), 
	.Q(cipher_sample[38]), 
	.D(FE_PHN1007_n359), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 cipher_sample_reg_46_ (.RN(reset_n), 
	.Q(cipher_sample[46]), 
	.D(FE_PHN3273_n351), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 cipher_sample_reg_54_ (.RN(reset_n), 
	.Q(cipher_sample[54]), 
	.D(FE_PHN1018_n343), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 cipher_sample_reg_62_ (.RN(reset_n), 
	.Q(cipher_sample[62]), 
	.D(FE_PHN941_n335), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 cipher_sample_reg_70_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[70]), 
	.D(FE_PHN1017_n327), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_78_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[78]), 
	.D(FE_PHN4854_n319), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_86_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[86]), 
	.D(FE_PHN832_n311), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_94_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[94]), 
	.D(FE_PHN3342_n303), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_102_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[102]), 
	.D(FE_PHN952_n295), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_110_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[110]), 
	.D(FE_PHN690_n287), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_118_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[118]), 
	.D(FE_PHN1335_n279), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 cipher_sample_reg_126_ (.RN(reset_n), 
	.Q(cipher_sample[126]), 
	.D(FE_PHN918_n271), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_5_ (.RN(reset_n), 
	.Q(cipher_sample[5]), 
	.D(FE_PHN1380_n392), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 cipher_sample_reg_13_ (.RN(reset_n), 
	.Q(cipher_sample[13]), 
	.D(FE_PHN851_n384), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_21_ (.RN(reset_n), 
	.Q(cipher_sample[21]), 
	.D(FE_PHN1030_n376), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 cipher_sample_reg_29_ (.RN(reset_n), 
	.Q(cipher_sample[29]), 
	.D(FE_PHN4962_n368), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_37_ (.RN(reset_n), 
	.Q(cipher_sample[37]), 
	.D(FE_PHN866_n360), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_45_ (.RN(reset_n), 
	.Q(cipher_sample[45]), 
	.D(FE_PHN725_n352), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_53_ (.RN(reset_n), 
	.Q(cipher_sample[53]), 
	.D(FE_PHN1360_n344), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_61_ (.RN(reset_n), 
	.Q(cipher_sample[61]), 
	.D(FE_PHN925_n336), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_69_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[69]), 
	.D(FE_PHN985_n328), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_77_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[77]), 
	.D(FE_PHN4666_n320), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_85_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[85]), 
	.D(FE_PHN826_n312), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_93_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[93]), 
	.D(FE_PHN729_n304), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_101_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[101]), 
	.D(FE_PHN1367_n296), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 cipher_sample_reg_109_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[109]), 
	.D(FE_PHN926_n288), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 cipher_sample_reg_117_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[117]), 
	.D(FE_PHN1028_n280), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 cipher_sample_reg_125_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[125]), 
	.D(FE_PHN2908_n272), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 cipher_sample_reg_4_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[4]), 
	.D(FE_PHN1261_n393), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 cipher_sample_reg_12_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[12]), 
	.D(FE_PHN842_n385), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_20_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[20]), 
	.D(FE_PHN1020_n377), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_28_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[28]), 
	.D(FE_PHN967_n369), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_36_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[36]), 
	.D(FE_PHN838_n361), 
	.CK(clk_48Mhz__L6_N44));
   DFFRHQX1 cipher_sample_reg_44_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[44]), 
	.D(FE_PHN3302_n353), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 cipher_sample_reg_52_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[52]), 
	.D(FE_PHN3327_n345), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 cipher_sample_reg_60_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[60]), 
	.D(FE_PHN1002_n337), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 cipher_sample_reg_68_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[68]), 
	.D(FE_PHN793_n329), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 cipher_sample_reg_76_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[76]), 
	.D(FE_PHN799_n321), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_84_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[84]), 
	.D(FE_PHN814_n313), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_92_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[92]), 
	.D(FE_PHN831_n305), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_100_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[100]), 
	.D(FE_PHN850_n297), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_108_ (.RN(FE_OFN53_reset_n), 
	.Q(cipher_sample[108]), 
	.D(FE_PHN801_n289), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_116_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[116]), 
	.D(FE_PHN978_n281), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 cipher_sample_reg_124_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_sample[124]), 
	.D(FE_PHN951_n273), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 cipher_sample_reg_3_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[3]), 
	.D(FE_PHN1107_n394), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_11_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[11]), 
	.D(FE_PHN761_n386), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_19_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[19]), 
	.D(FE_PHN778_n378), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 cipher_sample_reg_27_ (.RN(FE_OFN50_reset_n), 
	.Q(cipher_sample[27]), 
	.D(FE_PHN847_n370), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 cipher_sample_reg_35_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[35]), 
	.D(FE_PHN816_n362), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 cipher_sample_reg_43_ (.RN(FE_OFN50_reset_n), 
	.Q(cipher_sample[43]), 
	.D(FE_PHN804_n354), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 cipher_sample_reg_51_ (.RN(FE_OFN50_reset_n), 
	.Q(cipher_sample[51]), 
	.D(FE_PHN795_n346), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 cipher_sample_reg_59_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[59]), 
	.D(FE_PHN871_n338), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 cipher_sample_reg_67_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[67]), 
	.D(FE_PHN3308_n330), 
	.CK(clk_48Mhz__L6_N41));
   DFFRHQX1 cipher_sample_reg_75_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[75]), 
	.D(FE_PHN784_n322), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_83_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[83]), 
	.D(FE_PHN3330_n314), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_91_ (.RN(FE_OFN53_reset_n), 
	.Q(cipher_sample[91]), 
	.D(FE_PHN869_n306), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_99_ (.RN(FE_OFN53_reset_n), 
	.Q(cipher_sample[99]), 
	.D(FE_PHN839_n298), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_107_ (.RN(FE_OFN53_reset_n), 
	.Q(cipher_sample[107]), 
	.D(FE_PHN841_n290), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_115_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[115]), 
	.D(FE_PHN445_n282), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_123_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[123]), 
	.D(FE_PHN695_n274), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_2_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[2]), 
	.D(FE_PHN505_n395), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_10_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[10]), 
	.D(FE_PHN1289_n387), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_18_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[18]), 
	.D(FE_PHN858_n379), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_26_ (.RN(FE_OFN50_reset_n), 
	.Q(cipher_sample[26]), 
	.D(FE_PHN3335_n371), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_34_ (.RN(FE_OFN50_reset_n), 
	.Q(cipher_sample[34]), 
	.D(FE_PHN3378_n363), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_42_ (.RN(FE_OFN55_reset_n), 
	.Q(cipher_sample[42]), 
	.D(FE_PHN3388_n355), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_50_ (.RN(FE_OFN55_reset_n), 
	.Q(cipher_sample[50]), 
	.D(FE_PHN877_n347), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_58_ (.RN(FE_OFN55_reset_n), 
	.Q(cipher_sample[58]), 
	.D(FE_PHN859_n339), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_66_ (.RN(FE_OFN55_reset_n), 
	.Q(cipher_sample[66]), 
	.D(FE_PHN833_n331), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_74_ (.RN(FE_OFN39_reset_n), 
	.Q(cipher_sample[74]), 
	.D(FE_PHN3321_n323), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_82_ (.RN(FE_OFN39_reset_n), 
	.Q(cipher_sample[82]), 
	.D(FE_PHN636_n315), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_90_ (.RN(FE_OFN39_reset_n), 
	.Q(cipher_sample[90]), 
	.D(FE_PHN1299_n307), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_98_ (.RN(FE_OFN39_reset_n), 
	.Q(cipher_sample[98]), 
	.D(FE_PHN845_n299), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_106_ (.RN(FE_OFN39_reset_n), 
	.Q(cipher_sample[106]), 
	.D(FE_PHN629_n291), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_114_ (.RN(FE_OFN53_reset_n), 
	.Q(cipher_sample[114]), 
	.D(FE_PHN3365_n283), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_122_ (.RN(FE_OFN53_reset_n), 
	.Q(cipher_sample[122]), 
	.D(FE_PHN885_n275), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_1_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[1]), 
	.D(FE_PHN1172_n396), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_9_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[9]), 
	.D(FE_PHN863_n388), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_17_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[17]), 
	.D(FE_PHN787_n380), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_25_ (.RN(FE_OFN55_reset_n), 
	.Q(cipher_sample[25]), 
	.D(FE_PHN876_n372), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_33_ (.RN(FE_OFN55_reset_n), 
	.Q(cipher_sample[33]), 
	.D(FE_PHN693_n364), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_41_ (.RN(FE_OFN55_reset_n), 
	.Q(cipher_sample[41]), 
	.D(FE_PHN3341_n356), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_49_ (.RN(FE_OFN55_reset_n), 
	.Q(cipher_sample[49]), 
	.D(FE_PHN3289_n348), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_57_ (.RN(FE_OFN55_reset_n), 
	.Q(cipher_sample[57]), 
	.D(FE_PHN3322_n340), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_65_ (.RN(FE_OFN39_reset_n), 
	.Q(cipher_sample[65]), 
	.D(FE_PHN2990_n332), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_73_ (.RN(FE_OFN55_reset_n), 
	.Q(cipher_sample[73]), 
	.D(FE_PHN878_n324), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_81_ (.RN(FE_OFN55_reset_n), 
	.Q(cipher_sample[81]), 
	.D(FE_PHN3278_n316), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_89_ (.RN(FE_OFN39_reset_n), 
	.Q(cipher_sample[89]), 
	.D(FE_PHN790_n308), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_97_ (.RN(FE_OFN39_reset_n), 
	.Q(cipher_sample[97]), 
	.D(FE_PHN634_n300), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_105_ (.RN(FE_OFN53_reset_n), 
	.Q(cipher_sample[105]), 
	.D(FE_PHN1262_n292), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_113_ (.RN(FE_OFN53_reset_n), 
	.Q(cipher_sample[113]), 
	.D(FE_PHN759_n284), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_121_ (.RN(FE_OFN53_reset_n), 
	.Q(cipher_sample[121]), 
	.D(FE_PHN852_n276), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_0_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[0]), 
	.D(FE_PHN857_n397), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_8_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[8]), 
	.D(FE_PHN630_n389), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_16_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[16]), 
	.D(FE_PHN1288_n381), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_24_ (.RN(FE_OFN50_reset_n), 
	.Q(cipher_sample[24]), 
	.D(FE_PHN697_n373), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_32_ (.RN(FE_OFN55_reset_n), 
	.Q(cipher_sample[32]), 
	.D(FE_PHN1284_n365), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_40_ (.RN(FE_OFN55_reset_n), 
	.Q(cipher_sample[40]), 
	.D(FE_PHN781_n357), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_48_ (.RN(FE_OFN55_reset_n), 
	.Q(cipher_sample[48]), 
	.D(FE_PHN818_n349), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_56_ (.RN(FE_OFN55_reset_n), 
	.Q(cipher_sample[56]), 
	.D(FE_PHN868_n341), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_64_ (.RN(FE_OFN55_reset_n), 
	.Q(cipher_sample[64]), 
	.D(FE_PHN3260_n333), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_72_ (.RN(FE_OFN55_reset_n), 
	.Q(cipher_sample[72]), 
	.D(FE_PHN865_n325), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_80_ (.RN(FE_OFN39_reset_n), 
	.Q(cipher_sample[80]), 
	.D(FE_PHN809_n317), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_88_ (.RN(FE_OFN39_reset_n), 
	.Q(cipher_sample[88]), 
	.D(FE_PHN687_n309), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_96_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[96]), 
	.D(FE_PHN3252_n301), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_104_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[104]), 
	.D(FE_PHN358_n293), 
	.CK(clk_48Mhz__L6_N46));
   DFFRHQX1 cipher_sample_reg_112_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[112]), 
	.D(FE_PHN1265_n285), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 cipher_sample_reg_120_ (.RN(FE_OFN54_reset_n), 
	.Q(cipher_sample[120]), 
	.D(FE_PHN840_n277), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 rdy0_reg (.RN(FE_OFN53_reset_n), 
	.Q(rdy0), 
	.D(ready), 
	.CK(clk_48Mhz__L6_N47));
   DFFRHQX1 rdy2_reg (.RN(FE_OFN53_reset_n), 
	.Q(rdy2), 
	.D(FE_PHN5071_rdy1), 
	.CK(clk_48Mhz__L6_N43));
   DFFRHQX1 cipher_byte_reg_7_ (.RN(reset_n), 
	.Q(cipher_byte[7]), 
	.D(FE_PHN1449_n269), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 cipher_byte_reg_6_ (.RN(reset_n), 
	.Q(cipher_byte[6]), 
	.D(FE_PHN1419_n268), 
	.CK(clk_48Mhz__L6_N39));
   DFFRHQX1 cipher_byte_reg_5_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_byte[5]), 
	.D(FE_PHN1422_n267), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 cipher_byte_reg_4_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_byte[4]), 
	.D(FE_PHN1454_n266), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 cipher_byte_reg_3_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_byte[3]), 
	.D(FE_PHN1456_n265), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 cipher_byte_reg_2_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_byte[2]), 
	.D(FE_PHN1457_n264), 
	.CK(clk_48Mhz));
   DFFRHQX1 cipher_byte_reg_1_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_byte[1]), 
	.D(FE_PHN1458_n263), 
	.CK(clk_48Mhz));
   DFFRHQX1 cipher_byte_reg_0_ (.RN(FE_OFN46_reset_n), 
	.Q(cipher_byte[0]), 
	.D(FE_PHN2797_n262), 
	.CK(clk_48Mhz__L6_N45));
   DFFRHQX1 rdy1_reg (.RN(FE_OFN53_reset_n), 
	.Q(rdy1), 
	.D(FE_PHN5068_rdy0), 
	.CK(clk_48Mhz__L6_N47));
   AND2X2 U3 (.Y(n2), 
	.B(FE_OFN0_n1), 
	.A(n260));
   INVX1 U4 (.Y(n30), 
	.A(n2));
   INVX1 U5 (.Y(n28), 
	.A(n2));
   INVX1 U6 (.Y(n26), 
	.A(n2));
   INVX1 U7 (.Y(n25), 
	.A(n2));
   INVX1 U8 (.Y(n23), 
	.A(n2));
   INVX1 U13 (.Y(n4), 
	.A(n260));
   INVX1 U14 (.Y(n6), 
	.A(n260));
   INVX1 U15 (.Y(n7), 
	.A(n260));
   INVX1 U16 (.Y(n8), 
	.A(n260));
   INVX1 U17 (.Y(n10), 
	.A(n260));
   NAND3BX2 U34 (.Y(n1), 
	.C(FE_PHN124_rdy1), 
	.B(n54), 
	.AN(empty));
   OAI221XL U35 (.Y(n277), 
	.C0(n27), 
	.B1(n426), 
	.B0(n25), 
	.A1(FE_PHN1253_n425), 
	.A0(n1));
   NAND2X1 U36 (.Y(n27), 
	.B(n6), 
	.A(cipher_text[120]));
   OAI221XL U37 (.Y(n276), 
	.C0(n24), 
	.B1(n410), 
	.B0(n28), 
	.A1(FE_PHN3293_n409), 
	.A0(n1));
   NAND2X1 U38 (.Y(n24), 
	.B(n6), 
	.A(cipher_text[121]));
   OAI221XL U39 (.Y(n275), 
	.C0(n21), 
	.B1(n246), 
	.B0(n26), 
	.A1(n244), 
	.A0(n1));
   NAND2X1 U40 (.Y(n21), 
	.B(n6), 
	.A(cipher_text[122]));
   OAI221XL U41 (.Y(n274), 
	.C0(n18), 
	.B1(n214), 
	.B0(n23), 
	.A1(n212), 
	.A0(n1));
   NAND2X1 U42 (.Y(n18), 
	.B(n6), 
	.A(cipher_text[123]));
   OAI221XL U43 (.Y(n273), 
	.C0(n15), 
	.B1(n182), 
	.B0(n28), 
	.A1(FE_PHN3212_n180), 
	.A0(FE_OFN0_n1));
   NAND2X1 U44 (.Y(n15), 
	.B(n6), 
	.A(cipher_text[124]));
   OAI221XL U45 (.Y(n272), 
	.C0(n12), 
	.B1(n150), 
	.B0(n30), 
	.A1(FE_PHN3266_n148), 
	.A0(FE_OFN0_n1));
   NAND2X1 U46 (.Y(n12), 
	.B(n6), 
	.A(cipher_text[125]));
   OAI221XL U47 (.Y(n271), 
	.C0(n9), 
	.B1(n118), 
	.B0(n25), 
	.A1(n116), 
	.A0(FE_OFN0_n1));
   NAND2X1 U48 (.Y(n9), 
	.B(n6), 
	.A(cipher_text[126]));
   OAI221XL U49 (.Y(n270), 
	.C0(n5), 
	.B1(n86), 
	.B0(n30), 
	.A1(n84), 
	.A0(FE_OFN0_n1));
   NAND2X1 U50 (.Y(n5), 
	.B(n6), 
	.A(cipher_text[127]));
   OAI221XL U51 (.Y(n278), 
	.C0(n29), 
	.B1(n23), 
	.B0(n84), 
	.A1(n82), 
	.A0(FE_OFN0_n1));
   NAND2X1 U52 (.Y(n29), 
	.B(n6), 
	.A(cipher_text[119]));
   OAI221XL U53 (.Y(n285), 
	.C0(n43), 
	.B1(FE_PHN1253_n425), 
	.B0(n30), 
	.A1(FE_PHN3345_n424), 
	.A0(n1));
   NAND2X1 U54 (.Y(n43), 
	.B(n4), 
	.A(cipher_text[112]));
   OAI221XL U55 (.Y(n293), 
	.C0(n59), 
	.B1(FE_PHN3345_n424), 
	.B0(n28), 
	.A1(n423), 
	.A0(n1));
   NAND2X1 U56 (.Y(n59), 
	.B(n4), 
	.A(cipher_text[104]));
   OAI221XL U57 (.Y(n301), 
	.C0(n75), 
	.B1(n423), 
	.B0(n28), 
	.A1(n422), 
	.A0(n1));
   NAND2X1 U58 (.Y(n75), 
	.B(n6), 
	.A(cipher_text[96]));
   OAI221XL U59 (.Y(n309), 
	.C0(n91), 
	.B1(n422), 
	.B0(n26), 
	.A1(FE_PHN3246_n421), 
	.A0(n1));
   NAND2X1 U60 (.Y(n91), 
	.B(n7), 
	.A(cipher_text[88]));
   OAI221XL U61 (.Y(n317), 
	.C0(n107), 
	.B1(FE_PHN3246_n421), 
	.B0(n25), 
	.A1(FE_PHN2911_n420), 
	.A0(n1));
   NAND2X1 U62 (.Y(n107), 
	.B(n7), 
	.A(cipher_text[80]));
   OAI221XL U63 (.Y(n325), 
	.C0(n123), 
	.B1(FE_PHN2911_n420), 
	.B0(n25), 
	.A1(n419), 
	.A0(n1));
   NAND2X1 U64 (.Y(n123), 
	.B(n10), 
	.A(cipher_text[72]));
   OAI221XL U65 (.Y(n333), 
	.C0(n139), 
	.B1(n419), 
	.B0(n23), 
	.A1(FE_PHN3261_n418), 
	.A0(n1));
   NAND2X1 U66 (.Y(n139), 
	.B(n8), 
	.A(cipher_text[64]));
   OAI221XL U67 (.Y(n341), 
	.C0(n155), 
	.B1(FE_PHN3261_n418), 
	.B0(n23), 
	.A1(FE_PHN2910_n417), 
	.A0(n1));
   NAND2X1 U68 (.Y(n155), 
	.B(n8), 
	.A(cipher_text[56]));
   OAI221XL U69 (.Y(n349), 
	.C0(n171), 
	.B1(FE_PHN2910_n417), 
	.B0(n23), 
	.A1(n416), 
	.A0(n1));
   NAND2X1 U70 (.Y(n171), 
	.B(n10), 
	.A(cipher_text[48]));
   OAI221XL U71 (.Y(n357), 
	.C0(n187), 
	.B1(n416), 
	.B0(n25), 
	.A1(n415), 
	.A0(n1));
   NAND2X1 U72 (.Y(n187), 
	.B(n10), 
	.A(cipher_text[40]));
   OAI221XL U73 (.Y(n365), 
	.C0(n203), 
	.B1(n415), 
	.B0(n26), 
	.A1(FE_PHN3331_n414), 
	.A0(n1));
   NAND2X1 U74 (.Y(n203), 
	.B(n10), 
	.A(cipher_text[32]));
   OAI221XL U75 (.Y(n373), 
	.C0(n219), 
	.B1(FE_PHN3331_n414), 
	.B0(n26), 
	.A1(FE_PHN3255_n413), 
	.A0(n1));
   NAND2X1 U76 (.Y(n219), 
	.B(n8), 
	.A(cipher_text[24]));
   OAI221XL U77 (.Y(n381), 
	.C0(n235), 
	.B1(FE_PHN3255_n413), 
	.B0(n28), 
	.A1(n412), 
	.A0(n1));
   NAND2X1 U78 (.Y(n235), 
	.B(n7), 
	.A(cipher_text[16]));
   OAI221XL U79 (.Y(n389), 
	.C0(n251), 
	.B1(n412), 
	.B0(n30), 
	.A1(n411), 
	.A0(n1));
   NAND2X1 U80 (.Y(n251), 
	.B(n7), 
	.A(cipher_text[8]));
   OAI221XL U81 (.Y(n397), 
	.C0(n259), 
	.B1(n411), 
	.B0(n23), 
	.A1(n426), 
	.A0(n1));
   NAND2X1 U82 (.Y(n259), 
	.B(n6), 
	.A(cipher_text[0]));
   OAI221XL U83 (.Y(n284), 
	.C0(n41), 
	.B1(FE_PHN3293_n409), 
	.B0(n30), 
	.A1(FE_PHN3192_n408), 
	.A0(n1));
   NAND2X1 U84 (.Y(n41), 
	.B(n4), 
	.A(cipher_text[113]));
   OAI221XL U85 (.Y(n292), 
	.C0(n57), 
	.B1(FE_PHN3192_n408), 
	.B0(n28), 
	.A1(FE_PHN3329_n407), 
	.A0(n1));
   NAND2X1 U86 (.Y(n57), 
	.B(n4), 
	.A(cipher_text[105]));
   OAI221XL U87 (.Y(n300), 
	.C0(n73), 
	.B1(FE_PHN3329_n407), 
	.B0(n28), 
	.A1(FE_PHN3295_n406), 
	.A0(n1));
   NAND2X1 U88 (.Y(n73), 
	.B(n6), 
	.A(cipher_text[97]));
   OAI221XL U89 (.Y(n308), 
	.C0(n89), 
	.B1(FE_PHN3295_n406), 
	.B0(n26), 
	.A1(n405), 
	.A0(n1));
   NAND2X1 U90 (.Y(n89), 
	.B(n7), 
	.A(cipher_text[89]));
   OAI221XL U91 (.Y(n316), 
	.C0(n105), 
	.B1(n405), 
	.B0(n25), 
	.A1(n404), 
	.A0(n1));
   NAND2X1 U92 (.Y(n105), 
	.B(n7), 
	.A(cipher_text[81]));
   OAI221XL U93 (.Y(n324), 
	.C0(n121), 
	.B1(n404), 
	.B0(n25), 
	.A1(FE_PHN3362_n403), 
	.A0(n1));
   NAND2X1 U94 (.Y(n121), 
	.B(n8), 
	.A(cipher_text[73]));
   OAI221XL U95 (.Y(n332), 
	.C0(n137), 
	.B1(FE_PHN3362_n403), 
	.B0(n23), 
	.A1(n402), 
	.A0(n1));
   NAND2X1 U96 (.Y(n137), 
	.B(n8), 
	.A(cipher_text[65]));
   OAI221XL U97 (.Y(n340), 
	.C0(n153), 
	.B1(n402), 
	.B0(n23), 
	.A1(n401), 
	.A0(n1));
   NAND2X1 U98 (.Y(n153), 
	.B(n8), 
	.A(cipher_text[57]));
   OAI221XL U99 (.Y(n348), 
	.C0(n169), 
	.B1(n401), 
	.B0(n23), 
	.A1(n400), 
	.A0(n1));
   NAND2X1 U100 (.Y(n169), 
	.B(n10), 
	.A(cipher_text[49]));
   OAI221XL U101 (.Y(n356), 
	.C0(n185), 
	.B1(n400), 
	.B0(n25), 
	.A1(n399), 
	.A0(n1));
   NAND2X1 U102 (.Y(n185), 
	.B(n10), 
	.A(cipher_text[41]));
   OAI221XL U103 (.Y(n364), 
	.C0(n201), 
	.B1(n399), 
	.B0(n26), 
	.A1(n398), 
	.A0(n1));
   NAND2X1 U104 (.Y(n201), 
	.B(n10), 
	.A(cipher_text[33]));
   OAI221XL U105 (.Y(n372), 
	.C0(n217), 
	.B1(n398), 
	.B0(n26), 
	.A1(n261), 
	.A0(n1));
   NAND2X1 U106 (.Y(n217), 
	.B(n8), 
	.A(cipher_text[25]));
   OAI221XL U107 (.Y(n380), 
	.C0(n233), 
	.B1(n261), 
	.B0(n28), 
	.A1(FE_PHN2903_n250), 
	.A0(n1));
   NAND2X1 U108 (.Y(n233), 
	.B(n7), 
	.A(cipher_text[17]));
   OAI221XL U109 (.Y(n388), 
	.C0(n249), 
	.B1(FE_PHN2903_n250), 
	.B0(n30), 
	.A1(n248), 
	.A0(n1));
   NAND2X1 U110 (.Y(n249), 
	.B(n7), 
	.A(cipher_text[9]));
   OAI221XL U111 (.Y(n396), 
	.C0(n258), 
	.B1(n248), 
	.B0(n30), 
	.A1(n410), 
	.A0(n1));
   NAND2X1 U112 (.Y(n258), 
	.B(n7), 
	.A(cipher_text[1]));
   OAI221XL U113 (.Y(n283), 
	.C0(n39), 
	.B1(n244), 
	.B0(n30), 
	.A1(n242), 
	.A0(n1));
   NAND2X1 U114 (.Y(n39), 
	.B(n4), 
	.A(cipher_text[114]));
   OAI221XL U115 (.Y(n291), 
	.C0(n55), 
	.B1(n242), 
	.B0(n28), 
	.A1(FE_PHN2899_n240), 
	.A0(n1));
   NAND2X1 U116 (.Y(n55), 
	.B(n4), 
	.A(cipher_text[106]));
   OAI221XL U117 (.Y(n299), 
	.C0(n71), 
	.B1(FE_PHN2899_n240), 
	.B0(n28), 
	.A1(FE_PHN1255_n238), 
	.A0(n1));
   NAND2X1 U118 (.Y(n71), 
	.B(n6), 
	.A(cipher_text[98]));
   OAI221XL U119 (.Y(n307), 
	.C0(n87), 
	.B1(FE_PHN1255_n238), 
	.B0(n26), 
	.A1(n236), 
	.A0(n1));
   NAND2X1 U120 (.Y(n87), 
	.B(n7), 
	.A(cipher_text[90]));
   OAI221XL U121 (.Y(n315), 
	.C0(n103), 
	.B1(n236), 
	.B0(n25), 
	.A1(FE_PHN3267_n234), 
	.A0(n1));
   NAND2X1 U122 (.Y(n103), 
	.B(n7), 
	.A(cipher_text[82]));
   OAI221XL U123 (.Y(n323), 
	.C0(n119), 
	.B1(FE_PHN3267_n234), 
	.B0(n25), 
	.A1(n232), 
	.A0(n1));
   NAND2X1 U124 (.Y(n119), 
	.B(n4), 
	.A(cipher_text[74]));
   OAI221XL U125 (.Y(n331), 
	.C0(n135), 
	.B1(n232), 
	.B0(n23), 
	.A1(n230), 
	.A0(n1));
   NAND2X1 U126 (.Y(n135), 
	.B(n8), 
	.A(cipher_text[66]));
   OAI221XL U127 (.Y(n339), 
	.C0(n151), 
	.B1(n230), 
	.B0(n23), 
	.A1(FE_PHN3304_n228), 
	.A0(n1));
   NAND2X1 U128 (.Y(n151), 
	.B(n8), 
	.A(cipher_text[58]));
   OAI221XL U129 (.Y(n347), 
	.C0(n167), 
	.B1(FE_PHN3304_n228), 
	.B0(n23), 
	.A1(n226), 
	.A0(n1));
   NAND2X1 U130 (.Y(n167), 
	.B(n10), 
	.A(cipher_text[50]));
   OAI221XL U131 (.Y(n355), 
	.C0(n183), 
	.B1(n226), 
	.B0(n25), 
	.A1(n224), 
	.A0(n1));
   NAND2X1 U132 (.Y(n183), 
	.B(n10), 
	.A(cipher_text[42]));
   OAI221XL U133 (.Y(n363), 
	.C0(n199), 
	.B1(n224), 
	.B0(n26), 
	.A1(n222), 
	.A0(n1));
   NAND2X1 U134 (.Y(n199), 
	.B(n10), 
	.A(cipher_text[34]));
   OAI221XL U135 (.Y(n371), 
	.C0(n215), 
	.B1(n222), 
	.B0(n26), 
	.A1(FE_PHN2913_n220), 
	.A0(n1));
   NAND2X1 U136 (.Y(n215), 
	.B(n8), 
	.A(cipher_text[26]));
   OAI221XL U137 (.Y(n379), 
	.C0(n231), 
	.B1(FE_PHN2913_n220), 
	.B0(n28), 
	.A1(FE_PHN1259_n218), 
	.A0(n1));
   NAND2X1 U138 (.Y(n231), 
	.B(n7), 
	.A(cipher_text[18]));
   OAI221XL U139 (.Y(n387), 
	.C0(n247), 
	.B1(FE_PHN1259_n218), 
	.B0(n30), 
	.A1(n216), 
	.A0(n1));
   NAND2X1 U140 (.Y(n247), 
	.B(n7), 
	.A(cipher_text[10]));
   OAI221XL U141 (.Y(n395), 
	.C0(n257), 
	.B1(n216), 
	.B0(n30), 
	.A1(n246), 
	.A0(n1));
   NAND2X1 U142 (.Y(n257), 
	.B(n4), 
	.A(cipher_text[2]));
   OAI221XL U143 (.Y(n282), 
	.C0(n37), 
	.B1(n212), 
	.B0(n30), 
	.A1(n210), 
	.A0(n1));
   NAND2X1 U144 (.Y(n37), 
	.B(n4), 
	.A(cipher_text[115]));
   OAI221XL U145 (.Y(n290), 
	.C0(n53), 
	.B1(n210), 
	.B0(n30), 
	.A1(n208), 
	.A0(n1));
   NAND2X1 U146 (.Y(n53), 
	.B(n4), 
	.A(cipher_text[107]));
   OAI221XL U147 (.Y(n298), 
	.C0(n69), 
	.B1(n208), 
	.B0(n28), 
	.A1(n206), 
	.A0(n1));
   NAND2X1 U148 (.Y(n69), 
	.B(n6), 
	.A(cipher_text[99]));
   OAI221XL U149 (.Y(n306), 
	.C0(n85), 
	.B1(n206), 
	.B0(n26), 
	.A1(n204), 
	.A0(n1));
   NAND2X1 U150 (.Y(n85), 
	.B(n7), 
	.A(cipher_text[91]));
   OAI221XL U151 (.Y(n314), 
	.C0(n101), 
	.B1(n204), 
	.B0(n26), 
	.A1(n202), 
	.A0(n1));
   NAND2X1 U152 (.Y(n101), 
	.B(n7), 
	.A(cipher_text[83]));
   OAI221XL U153 (.Y(n322), 
	.C0(n117), 
	.B1(n202), 
	.B0(n25), 
	.A1(n200), 
	.A0(n1));
   NAND2X1 U154 (.Y(n117), 
	.B(n4), 
	.A(cipher_text[75]));
   OAI221XL U155 (.Y(n330), 
	.C0(n133), 
	.B1(n200), 
	.B0(n23), 
	.A1(n198), 
	.A0(n1));
   NAND2X1 U156 (.Y(n133), 
	.B(n8), 
	.A(cipher_text[67]));
   OAI221XL U157 (.Y(n338), 
	.C0(n149), 
	.B1(n198), 
	.B0(n23), 
	.A1(FE_PHN3356_n196), 
	.A0(n1));
   NAND2X1 U158 (.Y(n149), 
	.B(n8), 
	.A(cipher_text[59]));
   OAI221XL U159 (.Y(n346), 
	.C0(n165), 
	.B1(FE_PHN3356_n196), 
	.B0(n23), 
	.A1(FE_PHN3265_n194), 
	.A0(n1));
   NAND2X1 U160 (.Y(n165), 
	.B(n10), 
	.A(cipher_text[51]));
   OAI221XL U161 (.Y(n354), 
	.C0(n181), 
	.B1(FE_PHN3265_n194), 
	.B0(n25), 
	.A1(n192), 
	.A0(n1));
   NAND2X1 U162 (.Y(n181), 
	.B(n10), 
	.A(cipher_text[43]));
   OAI221XL U163 (.Y(n362), 
	.C0(n197), 
	.B1(n192), 
	.B0(n26), 
	.A1(n190), 
	.A0(n1));
   NAND2X1 U164 (.Y(n197), 
	.B(n10), 
	.A(cipher_text[35]));
   OAI221XL U165 (.Y(n370), 
	.C0(n213), 
	.B1(n190), 
	.B0(n26), 
	.A1(FE_PHN3263_n188), 
	.A0(n1));
   NAND2X1 U166 (.Y(n213), 
	.B(n8), 
	.A(cipher_text[27]));
   OAI221XL U167 (.Y(n378), 
	.C0(n229), 
	.B1(FE_PHN3263_n188), 
	.B0(n28), 
	.A1(FE_PHN3250_n186), 
	.A0(n1));
   NAND2X1 U168 (.Y(n229), 
	.B(n7), 
	.A(cipher_text[19]));
   OAI221XL U169 (.Y(n386), 
	.C0(n245), 
	.B1(FE_PHN3250_n186), 
	.B0(n30), 
	.A1(n184), 
	.A0(n1));
   NAND2X1 U170 (.Y(n245), 
	.B(n7), 
	.A(cipher_text[11]));
   OAI221XL U171 (.Y(n394), 
	.C0(n256), 
	.B1(n184), 
	.B0(n30), 
	.A1(n214), 
	.A0(n1));
   NAND2X1 U172 (.Y(n256), 
	.B(n4), 
	.A(cipher_text[3]));
   OAI221XL U173 (.Y(n281), 
	.C0(n35), 
	.B1(FE_PHN3212_n180), 
	.B0(n30), 
	.A1(n178), 
	.A0(FE_OFN0_n1));
   NAND2X1 U174 (.Y(n35), 
	.B(n6), 
	.A(cipher_text[116]));
   OAI221XL U175 (.Y(n289), 
	.C0(n51), 
	.B1(n178), 
	.B0(n30), 
	.A1(FE_PHN3241_n176), 
	.A0(n1));
   NAND2X1 U176 (.Y(n51), 
	.B(n4), 
	.A(cipher_text[108]));
   OAI221XL U177 (.Y(n297), 
	.C0(n67), 
	.B1(FE_PHN3241_n176), 
	.B0(n28), 
	.A1(n174), 
	.A0(n1));
   NAND2X1 U178 (.Y(n67), 
	.B(n6), 
	.A(cipher_text[100]));
   OAI221XL U179 (.Y(n305), 
	.C0(n83), 
	.B1(n174), 
	.B0(n26), 
	.A1(FE_PHN2904_n172), 
	.A0(n1));
   NAND2X1 U180 (.Y(n83), 
	.B(n6), 
	.A(cipher_text[92]));
   OAI221XL U181 (.Y(n313), 
	.C0(n99), 
	.B1(FE_PHN2904_n172), 
	.B0(n26), 
	.A1(n170), 
	.A0(n1));
   NAND2X1 U182 (.Y(n99), 
	.B(n7), 
	.A(cipher_text[84]));
   OAI221XL U183 (.Y(n321), 
	.C0(n115), 
	.B1(n170), 
	.B0(n25), 
	.A1(FE_PHN3269_n168), 
	.A0(n1));
   NAND2X1 U184 (.Y(n115), 
	.B(n4), 
	.A(cipher_text[76]));
   OAI221XL U185 (.Y(n329), 
	.C0(n131), 
	.B1(FE_PHN3269_n168), 
	.B0(n23), 
	.A1(n166), 
	.A0(n1));
   NAND2X1 U186 (.Y(n131), 
	.B(n4), 
	.A(cipher_text[68]));
   OAI221XL U187 (.Y(n337), 
	.C0(n147), 
	.B1(n166), 
	.B0(n23), 
	.A1(n164), 
	.A0(FE_OFN0_n1));
   NAND2X1 U188 (.Y(n147), 
	.B(n8), 
	.A(cipher_text[60]));
   OAI221XL U189 (.Y(n345), 
	.C0(n163), 
	.B1(n164), 
	.B0(n23), 
	.A1(n162), 
	.A0(FE_OFN0_n1));
   NAND2X1 U190 (.Y(n163), 
	.B(n10), 
	.A(cipher_text[52]));
   OAI221XL U191 (.Y(n353), 
	.C0(n179), 
	.B1(n162), 
	.B0(n25), 
	.A1(n160), 
	.A0(FE_OFN0_n1));
   NAND2X1 U192 (.Y(n179), 
	.B(n10), 
	.A(cipher_text[44]));
   OAI221XL U193 (.Y(n361), 
	.C0(n195), 
	.B1(n160), 
	.B0(n25), 
	.A1(n158), 
	.A0(FE_OFN0_n1));
   NAND2X1 U194 (.Y(n195), 
	.B(n10), 
	.A(cipher_text[36]));
   OAI221XL U195 (.Y(n369), 
	.C0(n211), 
	.B1(n158), 
	.B0(n26), 
	.A1(FE_PHN3220_n156), 
	.A0(FE_OFN0_n1));
   NAND2X1 U196 (.Y(n211), 
	.B(n8), 
	.A(cipher_text[28]));
   OAI221XL U197 (.Y(n377), 
	.C0(n227), 
	.B1(FE_PHN3220_n156), 
	.B0(n28), 
	.A1(n154), 
	.A0(FE_OFN0_n1));
   NAND2X1 U198 (.Y(n227), 
	.B(n8), 
	.A(cipher_text[20]));
   OAI221XL U199 (.Y(n385), 
	.C0(n243), 
	.B1(n154), 
	.B0(n28), 
	.A1(n152), 
	.A0(FE_OFN0_n1));
   NAND2X1 U200 (.Y(n243), 
	.B(n7), 
	.A(cipher_text[12]));
   OAI221XL U201 (.Y(n393), 
	.C0(n255), 
	.B1(n152), 
	.B0(n30), 
	.A1(n182), 
	.A0(FE_OFN0_n1));
   NAND2X1 U202 (.Y(n255), 
	.B(n4), 
	.A(cipher_text[4]));
   OAI221XL U203 (.Y(n280), 
	.C0(n33), 
	.B1(FE_PHN3266_n148), 
	.B0(n30), 
	.A1(n146), 
	.A0(FE_OFN0_n1));
   NAND2X1 U204 (.Y(n33), 
	.B(n6), 
	.A(cipher_text[117]));
   OAI221XL U205 (.Y(n288), 
	.C0(n49), 
	.B1(n146), 
	.B0(n30), 
	.A1(FE_PHN1237_n144), 
	.A0(FE_OFN0_n1));
   NAND2X1 U206 (.Y(n49), 
	.B(n4), 
	.A(cipher_text[109]));
   OAI221XL U207 (.Y(n296), 
	.C0(n65), 
	.B1(FE_PHN1237_n144), 
	.B0(n28), 
	.A1(n142), 
	.A0(FE_OFN0_n1));
   NAND2X1 U208 (.Y(n65), 
	.B(n6), 
	.A(cipher_text[101]));
   OAI221XL U209 (.Y(n304), 
	.C0(n81), 
	.B1(n142), 
	.B0(n26), 
	.A1(n140), 
	.A0(FE_OFN0_n1));
   NAND2X1 U210 (.Y(n81), 
	.B(n6), 
	.A(cipher_text[93]));
   OAI221XL U211 (.Y(n312), 
	.C0(n97), 
	.B1(n140), 
	.B0(n26), 
	.A1(FE_PHN2895_n138), 
	.A0(FE_OFN0_n1));
   NAND2X1 U212 (.Y(n97), 
	.B(n7), 
	.A(cipher_text[85]));
   OAI221XL U213 (.Y(n320), 
	.C0(n113), 
	.B1(FE_PHN2895_n138), 
	.B0(n25), 
	.A1(n136), 
	.A0(FE_OFN0_n1));
   NAND2X1 U214 (.Y(n113), 
	.B(n4), 
	.A(cipher_text[77]));
   OAI221XL U215 (.Y(n328), 
	.C0(n129), 
	.B1(n136), 
	.B0(n23), 
	.A1(n134), 
	.A0(FE_OFN0_n1));
   NAND2X1 U216 (.Y(n129), 
	.B(n8), 
	.A(cipher_text[69]));
   OAI221XL U217 (.Y(n336), 
	.C0(n145), 
	.B1(n134), 
	.B0(n23), 
	.A1(FE_PHN3202_n132), 
	.A0(FE_OFN0_n1));
   NAND2X1 U218 (.Y(n145), 
	.B(n8), 
	.A(cipher_text[61]));
   OAI221XL U219 (.Y(n344), 
	.C0(n161), 
	.B1(FE_PHN3202_n132), 
	.B0(n23), 
	.A1(FE_PHN3344_n130), 
	.A0(FE_OFN0_n1));
   NAND2X1 U220 (.Y(n161), 
	.B(n10), 
	.A(cipher_text[53]));
   OAI221XL U221 (.Y(n352), 
	.C0(n177), 
	.B1(FE_PHN3344_n130), 
	.B0(n25), 
	.A1(n128), 
	.A0(FE_OFN0_n1));
   NAND2X1 U222 (.Y(n177), 
	.B(n10), 
	.A(cipher_text[45]));
   OAI221XL U223 (.Y(n360), 
	.C0(n193), 
	.B1(n128), 
	.B0(n25), 
	.A1(n126), 
	.A0(FE_OFN0_n1));
   NAND2X1 U224 (.Y(n193), 
	.B(n10), 
	.A(cipher_text[37]));
   OAI221XL U225 (.Y(n368), 
	.C0(n209), 
	.B1(n126), 
	.B0(n26), 
	.A1(n124), 
	.A0(FE_OFN0_n1));
   NAND2X1 U226 (.Y(n209), 
	.B(n8), 
	.A(cipher_text[29]));
   OAI221XL U227 (.Y(n376), 
	.C0(n225), 
	.B1(n124), 
	.B0(n28), 
	.A1(n122), 
	.A0(FE_OFN0_n1));
   NAND2X1 U228 (.Y(n225), 
	.B(n8), 
	.A(cipher_text[21]));
   OAI221XL U229 (.Y(n384), 
	.C0(n241), 
	.B1(n122), 
	.B0(n28), 
	.A1(FE_PHN1258_n120), 
	.A0(FE_OFN0_n1));
   NAND2X1 U230 (.Y(n241), 
	.B(n7), 
	.A(cipher_text[13]));
   OAI221XL U231 (.Y(n392), 
	.C0(n254), 
	.B1(FE_PHN1258_n120), 
	.B0(n30), 
	.A1(n150), 
	.A0(FE_OFN0_n1));
   NAND2X1 U232 (.Y(n254), 
	.B(n4), 
	.A(cipher_text[5]));
   OAI221XL U233 (.Y(n279), 
	.C0(n31), 
	.B1(n116), 
	.B0(n30), 
	.A1(FE_PHN3259_n114), 
	.A0(FE_OFN0_n1));
   NAND2X1 U234 (.Y(n31), 
	.B(n6), 
	.A(cipher_text[118]));
   OAI221XL U235 (.Y(n287), 
	.C0(n47), 
	.B1(FE_PHN3259_n114), 
	.B0(n30), 
	.A1(n112), 
	.A0(FE_OFN0_n1));
   NAND2X1 U236 (.Y(n47), 
	.B(n4), 
	.A(cipher_text[110]));
   OAI221XL U237 (.Y(n295), 
	.C0(n63), 
	.B1(n112), 
	.B0(n28), 
	.A1(n110), 
	.A0(FE_OFN0_n1));
   NAND2X1 U238 (.Y(n63), 
	.B(n6), 
	.A(cipher_text[102]));
   OAI221XL U239 (.Y(n303), 
	.C0(n79), 
	.B1(n110), 
	.B0(n26), 
	.A1(n108), 
	.A0(FE_OFN0_n1));
   NAND2X1 U240 (.Y(n79), 
	.B(n6), 
	.A(cipher_text[94]));
   OAI221XL U241 (.Y(n311), 
	.C0(n95), 
	.B1(n108), 
	.B0(n26), 
	.A1(FE_PHN2909_n106), 
	.A0(FE_OFN0_n1));
   NAND2X1 U242 (.Y(n95), 
	.B(n7), 
	.A(cipher_text[86]));
   OAI221XL U243 (.Y(n319), 
	.C0(n111), 
	.B1(FE_PHN2909_n106), 
	.B0(n25), 
	.A1(n104), 
	.A0(FE_OFN0_n1));
   NAND2X1 U244 (.Y(n111), 
	.B(n7), 
	.A(cipher_text[78]));
   OAI221XL U245 (.Y(n327), 
	.C0(n127), 
	.B1(n104), 
	.B0(n23), 
	.A1(n102), 
	.A0(FE_OFN0_n1));
   NAND2X1 U246 (.Y(n127), 
	.B(n10), 
	.A(cipher_text[70]));
   OAI221XL U247 (.Y(n335), 
	.C0(n143), 
	.B1(n102), 
	.B0(n23), 
	.A1(FE_PHN3228_n100), 
	.A0(FE_OFN0_n1));
   NAND2X1 U248 (.Y(n143), 
	.B(n8), 
	.A(cipher_text[62]));
   OAI221XL U249 (.Y(n343), 
	.C0(n159), 
	.B1(FE_PHN3228_n100), 
	.B0(n23), 
	.A1(n98), 
	.A0(FE_OFN0_n1));
   NAND2X1 U250 (.Y(n159), 
	.B(n10), 
	.A(cipher_text[54]));
   OAI221XL U251 (.Y(n351), 
	.C0(n175), 
	.B1(n98), 
	.B0(n25), 
	.A1(FE_PHN3274_n96), 
	.A0(FE_OFN0_n1));
   NAND2X1 U252 (.Y(n175), 
	.B(n10), 
	.A(cipher_text[46]));
   OAI221XL U253 (.Y(n359), 
	.C0(n191), 
	.B1(FE_PHN3274_n96), 
	.B0(n25), 
	.A1(n94), 
	.A0(FE_OFN0_n1));
   NAND2X1 U254 (.Y(n191), 
	.B(n10), 
	.A(cipher_text[38]));
   OAI221XL U255 (.Y(n367), 
	.C0(n207), 
	.B1(n94), 
	.B0(n26), 
	.A1(n92), 
	.A0(FE_OFN0_n1));
   NAND2X1 U256 (.Y(n207), 
	.B(n8), 
	.A(cipher_text[30]));
   OAI221XL U257 (.Y(n375), 
	.C0(n223), 
	.B1(n92), 
	.B0(n28), 
	.A1(n90), 
	.A0(FE_OFN0_n1));
   NAND2X1 U258 (.Y(n223), 
	.B(n8), 
	.A(cipher_text[22]));
   OAI221XL U259 (.Y(n383), 
	.C0(n239), 
	.B1(n90), 
	.B0(n28), 
	.A1(FE_PHN1222_n88), 
	.A0(FE_OFN0_n1));
   NAND2X1 U260 (.Y(n239), 
	.B(n7), 
	.A(cipher_text[14]));
   OAI221XL U261 (.Y(n391), 
	.C0(n253), 
	.B1(FE_PHN1222_n88), 
	.B0(n30), 
	.A1(n118), 
	.A0(FE_OFN0_n1));
   NAND2X1 U262 (.Y(n253), 
	.B(n4), 
	.A(cipher_text[6]));
   OAI221XL U263 (.Y(n286), 
	.C0(n45), 
	.B1(n82), 
	.B0(n30), 
	.A1(n80), 
	.A0(FE_OFN0_n1));
   NAND2X1 U264 (.Y(n45), 
	.B(n4), 
	.A(cipher_text[111]));
   OAI221XL U265 (.Y(n294), 
	.C0(n61), 
	.B1(n80), 
	.B0(n28), 
	.A1(FE_PHN3271_n78), 
	.A0(FE_OFN0_n1));
   NAND2X1 U266 (.Y(n61), 
	.B(n6), 
	.A(cipher_text[103]));
   OAI221XL U267 (.Y(n302), 
	.C0(n77), 
	.B1(FE_PHN3271_n78), 
	.B0(n28), 
	.A1(FE_PHN3223_n76), 
	.A0(FE_OFN0_n1));
   NAND2X1 U268 (.Y(n77), 
	.B(n6), 
	.A(cipher_text[95]));
   OAI221XL U269 (.Y(n310), 
	.C0(n93), 
	.B1(FE_PHN3223_n76), 
	.B0(n26), 
	.A1(FE_PHN3256_n74), 
	.A0(FE_OFN0_n1));
   NAND2X1 U270 (.Y(n93), 
	.B(n7), 
	.A(cipher_text[87]));
   OAI221XL U271 (.Y(n318), 
	.C0(n109), 
	.B1(FE_PHN3256_n74), 
	.B0(n25), 
	.A1(n72), 
	.A0(FE_OFN0_n1));
   NAND2X1 U272 (.Y(n109), 
	.B(n4), 
	.A(cipher_text[79]));
   OAI221XL U273 (.Y(n326), 
	.C0(n125), 
	.B1(n72), 
	.B0(n25), 
	.A1(FE_PHN3225_n70), 
	.A0(FE_OFN0_n1));
   NAND2X1 U274 (.Y(n125), 
	.B(n6), 
	.A(cipher_text[71]));
   OAI221XL U275 (.Y(n334), 
	.C0(n141), 
	.B1(FE_PHN3225_n70), 
	.B0(n23), 
	.A1(FE_PHN3334_n68), 
	.A0(FE_OFN0_n1));
   NAND2X1 U276 (.Y(n141), 
	.B(n8), 
	.A(cipher_text[63]));
   OAI221XL U277 (.Y(n342), 
	.C0(n157), 
	.B1(FE_PHN3334_n68), 
	.B0(n23), 
	.A1(n66), 
	.A0(FE_OFN0_n1));
   NAND2X1 U278 (.Y(n157), 
	.B(n10), 
	.A(cipher_text[55]));
   OAI221XL U279 (.Y(n350), 
	.C0(n173), 
	.B1(n66), 
	.B0(n25), 
	.A1(FE_PHN3251_n64), 
	.A0(FE_OFN0_n1));
   NAND2X1 U280 (.Y(n173), 
	.B(n10), 
	.A(cipher_text[47]));
   OAI221XL U281 (.Y(n358), 
	.C0(n189), 
	.B1(FE_PHN3251_n64), 
	.B0(n25), 
	.A1(FE_PHN3314_n62), 
	.A0(FE_OFN0_n1));
   NAND2X1 U282 (.Y(n189), 
	.B(n10), 
	.A(cipher_text[39]));
   OAI221XL U283 (.Y(n366), 
	.C0(n205), 
	.B1(FE_PHN3314_n62), 
	.B0(n26), 
	.A1(n60), 
	.A0(FE_OFN0_n1));
   NAND2X1 U284 (.Y(n205), 
	.B(n8), 
	.A(cipher_text[31]));
   OAI221XL U285 (.Y(n374), 
	.C0(n221), 
	.B1(n60), 
	.B0(n28), 
	.A1(n58), 
	.A0(FE_OFN0_n1));
   NAND2X1 U286 (.Y(n221), 
	.B(n8), 
	.A(cipher_text[23]));
   OAI221XL U287 (.Y(n382), 
	.C0(n237), 
	.B1(n58), 
	.B0(n28), 
	.A1(FE_PHN1247_n56), 
	.A0(FE_OFN0_n1));
   NAND2X1 U288 (.Y(n237), 
	.B(n7), 
	.A(cipher_text[15]));
   OAI221XL U289 (.Y(n390), 
	.C0(n252), 
	.B1(FE_PHN1247_n56), 
	.B0(n30), 
	.A1(n86), 
	.A0(FE_OFN0_n1));
   NAND2X1 U290 (.Y(n252), 
	.B(n4), 
	.A(cipher_text[7]));
   NOR2BX1 U291 (.Y(cipher_byte_valid), 
	.B(FE_PHN124_rdy1), 
	.AN(rdy2));
   NAND3X1 U292 (.Y(n260), 
	.C(empty), 
	.B(n54), 
	.A(FE_PHN124_rdy1));
   OAI2BB2X1 U293 (.Y(n263), 
	.B1(n410), 
	.B0(FE_OFN0_n1), 
	.A1N(FE_OFN0_n1), 
	.A0N(cipher_byte[1]));
   OAI2BB2X1 U294 (.Y(n264), 
	.B1(n246), 
	.B0(FE_OFN0_n1), 
	.A1N(FE_OFN0_n1), 
	.A0N(cipher_byte[2]));
   OAI2BB2X1 U295 (.Y(n265), 
	.B1(n214), 
	.B0(FE_OFN0_n1), 
	.A1N(FE_OFN0_n1), 
	.A0N(cipher_byte[3]));
   OAI2BB2X1 U296 (.Y(n266), 
	.B1(n182), 
	.B0(FE_OFN0_n1), 
	.A1N(FE_OFN0_n1), 
	.A0N(cipher_byte[4]));
   OAI2BB2X1 U297 (.Y(n267), 
	.B1(n150), 
	.B0(FE_OFN0_n1), 
	.A1N(FE_OFN0_n1), 
	.A0N(cipher_byte[5]));
   OAI2BB2X1 U298 (.Y(n262), 
	.B1(n426), 
	.B0(FE_OFN0_n1), 
	.A1N(FE_OFN0_n1), 
	.A0N(cipher_byte[0]));
   OAI2BB2X1 U299 (.Y(n268), 
	.B1(n118), 
	.B0(FE_OFN0_n1), 
	.A1N(FE_OFN0_n1), 
	.A0N(cipher_byte[6]));
   OAI2BB2X1 U300 (.Y(n269), 
	.B1(n86), 
	.B0(FE_OFN0_n1), 
	.A1N(FE_OFN0_n1), 
	.A0N(cipher_byte[7]));
   INVX1 U301 (.Y(n54), 
	.A(FE_PHN115_rdy0));
   INVX1 U302 (.Y(n426), 
	.A(FE_PHN1455_cipher_sample_120_));
   INVX1 U303 (.Y(n410), 
	.A(cipher_sample[121]));
   INVX1 U304 (.Y(n246), 
	.A(FE_PHN3179_cipher_sample_122_));
   INVX1 U305 (.Y(n214), 
	.A(FE_PHN3177_cipher_sample_123_));
   INVX1 U306 (.Y(n182), 
	.A(FE_PHN2893_cipher_sample_124_));
   INVX1 U307 (.Y(n150), 
	.A(FE_PHN2891_cipher_sample_125_));
   INVX1 U308 (.Y(n118), 
	.A(FE_PHN2890_cipher_sample_126_));
   INVX1 U309 (.Y(n86), 
	.A(FE_PHN2892_cipher_sample_127_));
   INVX1 U310 (.Y(n84), 
	.A(FE_PHN3282_cipher_sample_119_));
   INVX1 U311 (.Y(n425), 
	.A(cipher_sample[112]));
   INVX1 U312 (.Y(n424), 
	.A(cipher_sample[104]));
   INVX1 U313 (.Y(n423), 
	.A(cipher_sample[96]));
   INVX1 U314 (.Y(n422), 
	.A(cipher_sample[88]));
   INVX1 U315 (.Y(n421), 
	.A(cipher_sample[80]));
   INVX1 U316 (.Y(n420), 
	.A(cipher_sample[72]));
   INVX1 U317 (.Y(n419), 
	.A(cipher_sample[64]));
   INVX1 U318 (.Y(n418), 
	.A(cipher_sample[56]));
   INVX1 U319 (.Y(n417), 
	.A(cipher_sample[48]));
   INVX1 U320 (.Y(n416), 
	.A(cipher_sample[40]));
   INVX1 U321 (.Y(n415), 
	.A(FE_PHN3244_cipher_sample_32_));
   INVX1 U322 (.Y(n414), 
	.A(cipher_sample[24]));
   INVX1 U323 (.Y(n413), 
	.A(cipher_sample[16]));
   INVX1 U324 (.Y(n412), 
	.A(FE_PHN3312_cipher_sample_8_));
   INVX1 U325 (.Y(n411), 
	.A(FE_PHN2898_cipher_sample_0_));
   INVX1 U326 (.Y(n409), 
	.A(cipher_sample[113]));
   INVX1 U327 (.Y(n408), 
	.A(cipher_sample[105]));
   INVX1 U328 (.Y(n407), 
	.A(cipher_sample[97]));
   INVX1 U329 (.Y(n406), 
	.A(cipher_sample[89]));
   INVX1 U330 (.Y(n405), 
	.A(cipher_sample[81]));
   INVX1 U331 (.Y(n404), 
	.A(FE_PHN3281_cipher_sample_73_));
   INVX1 U332 (.Y(n403), 
	.A(cipher_sample[65]));
   INVX1 U333 (.Y(n402), 
	.A(cipher_sample[57]));
   INVX1 U334 (.Y(n401), 
	.A(cipher_sample[49]));
   INVX1 U335 (.Y(n400), 
	.A(FE_PHN3290_cipher_sample_41_));
   INVX1 U336 (.Y(n399), 
	.A(cipher_sample[33]));
   INVX1 U337 (.Y(n398), 
	.A(FE_PHN2901_cipher_sample_25_));
   INVX1 U338 (.Y(n261), 
	.A(cipher_sample[17]));
   INVX1 U339 (.Y(n250), 
	.A(cipher_sample[9]));
   INVX1 U340 (.Y(n248), 
	.A(FE_PHN3360_cipher_sample_1_));
   INVX1 U341 (.Y(n244), 
	.A(FE_PHN2917_cipher_sample_114_));
   INVX1 U342 (.Y(n242), 
	.A(cipher_sample[106]));
   INVX1 U343 (.Y(n240), 
	.A(cipher_sample[98]));
   INVX1 U344 (.Y(n238), 
	.A(cipher_sample[90]));
   INVX1 U345 (.Y(n236), 
	.A(FE_PHN3371_cipher_sample_82_));
   INVX1 U346 (.Y(n234), 
	.A(cipher_sample[74]));
   INVX1 U347 (.Y(n232), 
	.A(cipher_sample[66]));
   INVX1 U348 (.Y(n230), 
	.A(FE_PHN3231_cipher_sample_58_));
   INVX1 U349 (.Y(n228), 
	.A(cipher_sample[50]));
   INVX1 U350 (.Y(n226), 
	.A(FE_PHN2919_cipher_sample_42_));
   INVX1 U351 (.Y(n224), 
	.A(cipher_sample[34]));
   INVX1 U352 (.Y(n222), 
	.A(cipher_sample[26]));
   INVX1 U353 (.Y(n220), 
	.A(cipher_sample[18]));
   INVX1 U354 (.Y(n218), 
	.A(cipher_sample[10]));
   INVX1 U355 (.Y(n216), 
	.A(FE_PHN2918_cipher_sample_2_));
   INVX1 U356 (.Y(n212), 
	.A(cipher_sample[115]));
   INVX1 U357 (.Y(n210), 
	.A(FE_PHN3238_cipher_sample_107_));
   INVX1 U358 (.Y(n208), 
	.A(cipher_sample[99]));
   INVX1 U359 (.Y(n206), 
	.A(FE_PHN3233_cipher_sample_91_));
   INVX1 U360 (.Y(n204), 
	.A(cipher_sample[83]));
   INVX1 U361 (.Y(n202), 
	.A(cipher_sample[75]));
   INVX1 U362 (.Y(n200), 
	.A(FE_PHN3217_cipher_sample_67_));
   INVX1 U363 (.Y(n198), 
	.A(FE_PHN3309_cipher_sample_59_));
   INVX1 U364 (.Y(n196), 
	.A(cipher_sample[51]));
   INVX1 U365 (.Y(n194), 
	.A(cipher_sample[43]));
   INVX1 U366 (.Y(n192), 
	.A(FE_PHN3325_cipher_sample_35_));
   INVX1 U367 (.Y(n190), 
	.A(cipher_sample[27]));
   INVX1 U368 (.Y(n188), 
	.A(cipher_sample[19]));
   INVX1 U369 (.Y(n186), 
	.A(cipher_sample[11]));
   INVX1 U370 (.Y(n184), 
	.A(FE_PHN2897_cipher_sample_3_));
   INVX1 U371 (.Y(n180), 
	.A(cipher_sample[116]));
   INVX1 U372 (.Y(n178), 
	.A(cipher_sample[108]));
   INVX1 U373 (.Y(n176), 
	.A(cipher_sample[100]));
   INVX1 U374 (.Y(n174), 
	.A(cipher_sample[92]));
   INVX1 U375 (.Y(n172), 
	.A(cipher_sample[84]));
   INVX1 U376 (.Y(n170), 
	.A(cipher_sample[76]));
   INVX1 U377 (.Y(n168), 
	.A(cipher_sample[68]));
   INVX1 U378 (.Y(n166), 
	.A(FE_PHN3277_cipher_sample_60_));
   INVX1 U379 (.Y(n164), 
	.A(FE_PHN3296_cipher_sample_52_));
   INVX1 U380 (.Y(n162), 
	.A(cipher_sample[44]));
   INVX1 U381 (.Y(n160), 
	.A(FE_PHN3301_cipher_sample_36_));
   INVX1 U382 (.Y(n158), 
	.A(cipher_sample[28]));
   INVX1 U383 (.Y(n156), 
	.A(cipher_sample[20]));
   INVX1 U384 (.Y(n154), 
	.A(FE_PHN2915_cipher_sample_12_));
   INVX1 U385 (.Y(n152), 
	.A(FE_PHN1254_cipher_sample_4_));
   INVX1 U386 (.Y(n148), 
	.A(cipher_sample[117]));
   INVX1 U387 (.Y(n146), 
	.A(FE_PHN2914_cipher_sample_109_));
   INVX1 U388 (.Y(n144), 
	.A(cipher_sample[101]));
   INVX1 U389 (.Y(n142), 
	.A(FE_PHN3351_cipher_sample_93_));
   INVX1 U390 (.Y(n140), 
	.A(cipher_sample[85]));
   INVX1 U391 (.Y(n138), 
	.A(cipher_sample[77]));
   INVX1 U392 (.Y(n136), 
	.A(cipher_sample[69]));
   INVX1 U393 (.Y(n134), 
	.A(cipher_sample[61]));
   INVX1 U394 (.Y(n132), 
	.A(cipher_sample[53]));
   INVX1 U395 (.Y(n130), 
	.A(cipher_sample[45]));
   INVX1 U396 (.Y(n128), 
	.A(FE_PHN2907_cipher_sample_37_));
   INVX1 U397 (.Y(n126), 
	.A(cipher_sample[29]));
   INVX1 U398 (.Y(n124), 
	.A(FE_PHN2912_cipher_sample_21_));
   INVX1 U399 (.Y(n122), 
	.A(FE_PHN3340_cipher_sample_13_));
   INVX1 U400 (.Y(n120), 
	.A(cipher_sample[5]));
   INVX1 U401 (.Y(n116), 
	.A(FE_PHN3191_cipher_sample_118_));
   INVX1 U402 (.Y(n114), 
	.A(cipher_sample[110]));
   INVX1 U403 (.Y(n112), 
	.A(FE_PHN3216_cipher_sample_102_));
   INVX1 U404 (.Y(n110), 
	.A(FE_PHN2902_cipher_sample_94_));
   INVX1 U405 (.Y(n108), 
	.A(cipher_sample[86]));
   INVX1 U406 (.Y(n106), 
	.A(cipher_sample[78]));
   INVX1 U407 (.Y(n104), 
	.A(cipher_sample[70]));
   INVX1 U408 (.Y(n102), 
	.A(cipher_sample[62]));
   INVX1 U409 (.Y(n100), 
	.A(cipher_sample[54]));
   INVX1 U410 (.Y(n98), 
	.A(cipher_sample[46]));
   INVX1 U411 (.Y(n96), 
	.A(cipher_sample[38]));
   INVX1 U412 (.Y(n94), 
	.A(FE_PHN3326_cipher_sample_30_));
   INVX1 U413 (.Y(n92), 
	.A(FE_PHN2906_cipher_sample_22_));
   INVX1 U414 (.Y(n90), 
	.A(FE_PHN3353_cipher_sample_14_));
   INVX1 U415 (.Y(n88), 
	.A(cipher_sample[6]));
   INVX1 U416 (.Y(n82), 
	.A(FE_PHN2896_cipher_sample_111_));
   INVX1 U417 (.Y(n80), 
	.A(cipher_sample[103]));
   INVX1 U418 (.Y(n78), 
	.A(cipher_sample[95]));
   INVX1 U419 (.Y(n76), 
	.A(cipher_sample[87]));
   INVX1 U420 (.Y(n74), 
	.A(cipher_sample[79]));
   INVX1 U421 (.Y(n72), 
	.A(cipher_sample[71]));
   INVX1 U422 (.Y(n70), 
	.A(cipher_sample[63]));
   INVX1 U423 (.Y(n68), 
	.A(cipher_sample[55]));
   INVX1 U424 (.Y(n66), 
	.A(cipher_sample[47]));
   INVX1 U425 (.Y(n64), 
	.A(cipher_sample[39]));
   INVX1 U426 (.Y(n62), 
	.A(cipher_sample[31]));
   INVX1 U427 (.Y(n60), 
	.A(FE_PHN3316_cipher_sample_23_));
   INVX1 U428 (.Y(n58), 
	.A(FE_PHN2916_cipher_sample_15_));
   INVX1 U429 (.Y(n56), 
	.A(cipher_sample[7]));
endmodule

module aes_top (
	reset_p, 
	clk_48Mhz, 
	plain_byte_in, 
	plain_byte_valid, 
	plain_finish, 
	empty, 
	cipher_byte_out, 
	cipher_byte_valid, 
	trig);
   input reset_p;
   input clk_48Mhz;
   input [7:0] plain_byte_in;
   input plain_byte_valid;
   input plain_finish;
   input empty;
   output [7:0] cipher_byte_out;
   output cipher_byte_valid;
   output trig;

   // Internal wires
   wire FE_PHN5173_reset_n;
   wire FE_PHN2803_reset_n;
   wire FE_PHN110_reset_n;
   wire clk_48Mhz__L6_N47;
   wire clk_48Mhz__L6_N46;
   wire clk_48Mhz__L6_N45;
   wire clk_48Mhz__L6_N44;
   wire clk_48Mhz__L6_N43;
   wire clk_48Mhz__L6_N42;
   wire clk_48Mhz__L6_N41;
   wire clk_48Mhz__L6_N40;
   wire clk_48Mhz__L6_N39;
   wire clk_48Mhz__L6_N38;
   wire clk_48Mhz__L6_N37;
   wire clk_48Mhz__L6_N36;
   wire clk_48Mhz__L6_N35;
   wire clk_48Mhz__L6_N34;
   wire clk_48Mhz__L6_N33;
   wire clk_48Mhz__L6_N32;
   wire clk_48Mhz__L6_N31;
   wire clk_48Mhz__L6_N30;
   wire clk_48Mhz__L6_N29;
   wire clk_48Mhz__L6_N28;
   wire clk_48Mhz__L6_N27;
   wire clk_48Mhz__L6_N26;
   wire clk_48Mhz__L6_N25;
   wire clk_48Mhz__L6_N24;
   wire clk_48Mhz__L6_N23;
   wire clk_48Mhz__L6_N22;
   wire clk_48Mhz__L6_N21;
   wire clk_48Mhz__L6_N20;
   wire clk_48Mhz__L6_N19;
   wire clk_48Mhz__L6_N18;
   wire clk_48Mhz__L6_N17;
   wire clk_48Mhz__L6_N16;
   wire clk_48Mhz__L6_N15;
   wire clk_48Mhz__L6_N14;
   wire clk_48Mhz__L6_N13;
   wire clk_48Mhz__L6_N12;
   wire clk_48Mhz__L6_N11;
   wire clk_48Mhz__L6_N10;
   wire clk_48Mhz__L6_N9;
   wire clk_48Mhz__L6_N8;
   wire clk_48Mhz__L6_N7;
   wire clk_48Mhz__L6_N6;
   wire clk_48Mhz__L6_N5;
   wire clk_48Mhz__L6_N4;
   wire clk_48Mhz__L6_N3;
   wire clk_48Mhz__L6_N2;
   wire clk_48Mhz__L6_N1;
   wire clk_48Mhz__L6_N0;
   wire clk_48Mhz__L5_N0;
   wire clk_48Mhz__L4_N0;
   wire clk_48Mhz__L3_N0;
   wire clk_48Mhz__L2_N0;
   wire clk_48Mhz__L1_N0;
   wire FE_OFN58_reset_n;
   wire FE_OFN56_reset_n;
   wire FE_OFN55_reset_n;
   wire FE_OFN54_reset_n;
   wire FE_OFN53_reset_n;
   wire FE_OFN51_reset_n;
   wire FE_OFN50_reset_n;
   wire FE_OFN49_reset_n;
   wire FE_OFN48_reset_n;
   wire FE_OFN47_reset_n;
   wire FE_OFN46_reset_n;
   wire FE_OFN45_reset_n;
   wire FE_OFN44_reset_n;
   wire FE_OFN43_reset_n;
   wire FE_OFN42_reset_n;
   wire FE_OFN40_reset_n;
   wire FE_OFN39_reset_n;
   wire FE_OFN38_reset_n;
   wire FE_OFN37_reset_n;
   wire FE_OFN34_reset_n;
   wire reset_n;
   wire init;
   wire next;
   wire ready;
   wire [255:0] Din;
   wire [127:0] Dout;

   DLY2X1 FE_PHC5173_reset_n (.Y(FE_PHN5173_reset_n), 
	.A(reset_n));
   DLY4X1 FE_PHC2803_reset_n (.Y(FE_PHN2803_reset_n), 
	.A(FE_PHN110_reset_n));
   DLY4X1 FE_PHC110_reset_n (.Y(FE_PHN110_reset_n), 
	.A(FE_PHN5173_reset_n));
   CLKBUFX8 clk_48Mhz__L6_I47 (.Y(clk_48Mhz__L6_N47), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I46 (.Y(clk_48Mhz__L6_N46), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I45 (.Y(clk_48Mhz__L6_N45), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I44 (.Y(clk_48Mhz__L6_N44), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I43 (.Y(clk_48Mhz__L6_N43), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I42 (.Y(clk_48Mhz__L6_N42), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I41 (.Y(clk_48Mhz__L6_N41), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I40 (.Y(clk_48Mhz__L6_N40), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I39 (.Y(clk_48Mhz__L6_N39), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I38 (.Y(clk_48Mhz__L6_N38), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I37 (.Y(clk_48Mhz__L6_N37), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I36 (.Y(clk_48Mhz__L6_N36), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I35 (.Y(clk_48Mhz__L6_N35), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I34 (.Y(clk_48Mhz__L6_N34), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I33 (.Y(clk_48Mhz__L6_N33), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I32 (.Y(clk_48Mhz__L6_N32), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I31 (.Y(clk_48Mhz__L6_N31), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I30 (.Y(clk_48Mhz__L6_N30), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I29 (.Y(clk_48Mhz__L6_N29), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I28 (.Y(clk_48Mhz__L6_N28), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I27 (.Y(clk_48Mhz__L6_N27), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I26 (.Y(clk_48Mhz__L6_N26), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I25 (.Y(clk_48Mhz__L6_N25), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I24 (.Y(clk_48Mhz__L6_N24), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I23 (.Y(clk_48Mhz__L6_N23), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I22 (.Y(clk_48Mhz__L6_N22), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I21 (.Y(clk_48Mhz__L6_N21), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I20 (.Y(clk_48Mhz__L6_N20), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I19 (.Y(clk_48Mhz__L6_N19), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I18 (.Y(clk_48Mhz__L6_N18), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I17 (.Y(clk_48Mhz__L6_N17), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I16 (.Y(clk_48Mhz__L6_N16), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I15 (.Y(clk_48Mhz__L6_N15), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I14 (.Y(clk_48Mhz__L6_N14), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I13 (.Y(clk_48Mhz__L6_N13), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I12 (.Y(clk_48Mhz__L6_N12), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I11 (.Y(clk_48Mhz__L6_N11), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I10 (.Y(clk_48Mhz__L6_N10), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I9 (.Y(clk_48Mhz__L6_N9), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I8 (.Y(clk_48Mhz__L6_N8), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I7 (.Y(clk_48Mhz__L6_N7), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I6 (.Y(clk_48Mhz__L6_N6), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I5 (.Y(clk_48Mhz__L6_N5), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I4 (.Y(clk_48Mhz__L6_N4), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I3 (.Y(clk_48Mhz__L6_N3), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I2 (.Y(clk_48Mhz__L6_N2), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I1 (.Y(clk_48Mhz__L6_N1), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX8 clk_48Mhz__L6_I0 (.Y(clk_48Mhz__L6_N0), 
	.A(clk_48Mhz__L5_N0));
   CLKBUFX20 clk_48Mhz__L5_I0 (.Y(clk_48Mhz__L5_N0), 
	.A(clk_48Mhz__L4_N0));
   CLKBUFX4 clk_48Mhz__L4_I0 (.Y(clk_48Mhz__L4_N0), 
	.A(clk_48Mhz__L3_N0));
   CLKBUFX4 clk_48Mhz__L3_I0 (.Y(clk_48Mhz__L3_N0), 
	.A(clk_48Mhz__L2_N0));
   CLKBUFX4 clk_48Mhz__L2_I0 (.Y(clk_48Mhz__L2_N0), 
	.A(clk_48Mhz__L1_N0));
   CLKBUFX20 clk_48Mhz__L1_I0 (.Y(clk_48Mhz__L1_N0), 
	.A(clk_48Mhz));
   CLKINVX3 FE_OFC58_reset_n (.Y(FE_OFN58_reset_n), 
	.A(FE_OFN48_reset_n));
   INVX1 FE_OFC56_reset_n (.Y(FE_OFN56_reset_n), 
	.A(FE_OFN48_reset_n));
   CLKINVX2 FE_OFC55_reset_n (.Y(FE_OFN55_reset_n), 
	.A(FE_OFN48_reset_n));
   CLKBUFX2 FE_OFC54_reset_n (.Y(FE_OFN54_reset_n), 
	.A(FE_OFN50_reset_n));
   CLKBUFX3 FE_OFC53_reset_n (.Y(FE_OFN53_reset_n), 
	.A(FE_OFN46_reset_n));
   CLKBUFX2 FE_OFC51_reset_n (.Y(FE_OFN51_reset_n), 
	.A(FE_OFN38_reset_n));
   CLKBUFX2 FE_OFC50_reset_n (.Y(FE_OFN50_reset_n), 
	.A(FE_OFN38_reset_n));
   CLKBUFX2 FE_OFC49_reset_n (.Y(FE_OFN49_reset_n), 
	.A(FE_OFN40_reset_n));
   INVX1 FE_OFC48_reset_n (.Y(FE_OFN48_reset_n), 
	.A(FE_OFN43_reset_n));
   CLKBUFX2 FE_OFC47_reset_n (.Y(FE_OFN47_reset_n), 
	.A(FE_OFN40_reset_n));
   CLKBUFX3 FE_OFC46_reset_n (.Y(FE_OFN46_reset_n), 
	.A(FE_OFN39_reset_n));
   CLKBUFX2 FE_OFC45_reset_n (.Y(FE_OFN45_reset_n), 
	.A(FE_OFN37_reset_n));
   CLKINVX3 FE_OFC44_reset_n (.Y(FE_OFN44_reset_n), 
	.A(FE_OFN34_reset_n));
   CLKINVX2 FE_OFC43_reset_n (.Y(FE_OFN43_reset_n), 
	.A(FE_OFN34_reset_n));
   CLKINVX3 FE_OFC42_reset_n (.Y(FE_OFN42_reset_n), 
	.A(FE_OFN34_reset_n));
   CLKINVX2 FE_OFC40_reset_n (.Y(FE_OFN40_reset_n), 
	.A(FE_OFN34_reset_n));
   CLKINVX2 FE_OFC39_reset_n (.Y(FE_OFN39_reset_n), 
	.A(FE_OFN34_reset_n));
   CLKINVX3 FE_OFC38_reset_n (.Y(FE_OFN38_reset_n), 
	.A(FE_OFN34_reset_n));
   CLKINVX3 FE_OFC37_reset_n (.Y(FE_OFN37_reset_n), 
	.A(FE_OFN34_reset_n));
   INVX2 FE_OFC34_reset_n (.Y(FE_OFN34_reset_n), 
	.A(FE_PHN2803_reset_n));
   INVX1 U1 (.Y(reset_n), 
	.A(reset_p));
   control control (.clk(clk_48Mhz__L6_N18), 
	.rst_n(FE_OFN53_reset_n), 
	.init(init), 
	.next(next), 
	.trig(trig), 
	.clk_48Mhz__L6_N43(clk_48Mhz__L6_N43));
   aes_core aes_core (.clk(clk_48Mhz__L6_N0), 
	.reset_n(FE_OFN34_reset_n), 
	.init(init), 
	.next(next), 
	.ready(ready), 
	.key({ Din[255],
		Din[254],
		Din[253],
		Din[252],
		Din[251],
		Din[250],
		Din[249],
		Din[248],
		Din[247],
		Din[246],
		Din[245],
		Din[244],
		Din[243],
		Din[242],
		Din[241],
		Din[240],
		Din[239],
		Din[238],
		Din[237],
		Din[236],
		Din[235],
		Din[234],
		Din[233],
		Din[232],
		Din[231],
		Din[230],
		Din[229],
		Din[228],
		Din[227],
		Din[226],
		Din[225],
		Din[224],
		Din[223],
		Din[222],
		Din[221],
		Din[220],
		Din[219],
		Din[218],
		Din[217],
		Din[216],
		Din[215],
		Din[214],
		Din[213],
		Din[212],
		Din[211],
		Din[210],
		Din[209],
		Din[208],
		Din[207],
		Din[206],
		Din[205],
		Din[204],
		Din[203],
		Din[202],
		Din[201],
		Din[200],
		Din[199],
		Din[198],
		Din[197],
		Din[196],
		Din[195],
		Din[194],
		Din[193],
		Din[192],
		Din[191],
		Din[190],
		Din[189],
		Din[188],
		Din[187],
		Din[186],
		Din[185],
		Din[184],
		Din[183],
		Din[182],
		Din[181],
		Din[180],
		Din[179],
		Din[178],
		Din[177],
		Din[176],
		Din[175],
		Din[174],
		Din[173],
		Din[172],
		Din[171],
		Din[170],
		Din[169],
		Din[168],
		Din[167],
		Din[166],
		Din[165],
		Din[164],
		Din[163],
		Din[162],
		Din[161],
		Din[160],
		Din[159],
		Din[158],
		Din[157],
		Din[156],
		Din[155],
		Din[154],
		Din[153],
		Din[152],
		Din[151],
		Din[150],
		Din[149],
		Din[148],
		Din[147],
		Din[146],
		Din[145],
		Din[144],
		Din[143],
		Din[142],
		Din[141],
		Din[140],
		Din[139],
		Din[138],
		Din[137],
		Din[136],
		Din[135],
		Din[134],
		Din[133],
		Din[132],
		Din[131],
		Din[130],
		Din[129],
		Din[128] }), 
	.block({ Din[127],
		Din[126],
		Din[125],
		Din[124],
		Din[123],
		Din[122],
		Din[121],
		Din[120],
		Din[119],
		Din[118],
		Din[117],
		Din[116],
		Din[115],
		Din[114],
		Din[113],
		Din[112],
		Din[111],
		Din[110],
		Din[109],
		Din[108],
		Din[107],
		Din[106],
		Din[105],
		Din[104],
		Din[103],
		Din[102],
		Din[101],
		Din[100],
		Din[99],
		Din[98],
		Din[97],
		Din[96],
		Din[95],
		Din[94],
		Din[93],
		Din[92],
		Din[91],
		Din[90],
		Din[89],
		Din[88],
		Din[87],
		Din[86],
		Din[85],
		Din[84],
		Din[83],
		Din[82],
		Din[81],
		Din[80],
		Din[79],
		Din[78],
		Din[77],
		Din[76],
		Din[75],
		Din[74],
		Din[73],
		Din[72],
		Din[71],
		Din[70],
		Din[69],
		Din[68],
		Din[67],
		Din[66],
		Din[65],
		Din[64],
		Din[63],
		Din[62],
		Din[61],
		Din[60],
		Din[59],
		Din[58],
		Din[57],
		Din[56],
		Din[55],
		Din[54],
		Din[53],
		Din[52],
		Din[51],
		Din[50],
		Din[49],
		Din[48],
		Din[47],
		Din[46],
		Din[45],
		Din[44],
		Din[43],
		Din[42],
		Din[41],
		Din[40],
		Din[39],
		Din[38],
		Din[37],
		Din[36],
		Din[35],
		Din[34],
		Din[33],
		Din[32],
		Din[31],
		Din[30],
		Din[29],
		Din[28],
		Din[27],
		Din[26],
		Din[25],
		Din[24],
		Din[23],
		Din[22],
		Din[21],
		Din[20],
		Din[19],
		Din[18],
		Din[17],
		Din[16],
		Din[15],
		Din[14],
		Din[13],
		Din[12],
		Din[11],
		Din[10],
		Din[9],
		Din[8],
		Din[7],
		Din[6],
		Din[5],
		Din[4],
		Din[3],
		Din[2],
		Din[1],
		Din[0] }), 
	.result(Dout), 
	.FE_OFN37_reset_n(FE_OFN37_reset_n), 
	.FE_OFN38_reset_n(FE_OFN38_reset_n), 
	.FE_OFN39_reset_n(FE_OFN39_reset_n), 
	.FE_OFN40_reset_n(FE_OFN40_reset_n), 
	.FE_OFN42_reset_n(FE_OFN42_reset_n), 
	.FE_OFN43_reset_n(FE_OFN43_reset_n), 
	.FE_OFN44_reset_n(FE_OFN44_reset_n), 
	.FE_OFN45_reset_n(FE_OFN45_reset_n), 
	.FE_OFN46_reset_n(FE_OFN46_reset_n), 
	.FE_OFN47_reset_n(FE_OFN47_reset_n), 
	.FE_OFN48_reset_n(FE_OFN48_reset_n), 
	.FE_OFN49_reset_n(FE_OFN49_reset_n), 
	.FE_OFN50_reset_n(FE_OFN50_reset_n), 
	.FE_OFN51_reset_n(FE_OFN51_reset_n), 
	.FE_OFN53_reset_n(FE_OFN53_reset_n), 
	.FE_OFN54_reset_n(FE_OFN54_reset_n), 
	.FE_OFN55_reset_n(FE_OFN55_reset_n), 
	.FE_OFN56_reset_n(FE_OFN56_reset_n), 
	.FE_OFN58_reset_n(FE_OFN58_reset_n), 
	.clk_48Mhz__L6_N1(clk_48Mhz__L6_N1), 
	.clk_48Mhz__L6_N10(clk_48Mhz__L6_N10), 
	.clk_48Mhz__L6_N11(clk_48Mhz__L6_N11), 
	.clk_48Mhz__L6_N12(clk_48Mhz__L6_N12), 
	.clk_48Mhz__L6_N13(clk_48Mhz__L6_N13), 
	.clk_48Mhz__L6_N14(clk_48Mhz__L6_N14), 
	.clk_48Mhz__L6_N15(clk_48Mhz__L6_N15), 
	.clk_48Mhz__L6_N16(clk_48Mhz__L6_N16), 
	.clk_48Mhz__L6_N17(clk_48Mhz__L6_N17), 
	.clk_48Mhz__L6_N18(clk_48Mhz__L6_N18), 
	.clk_48Mhz__L6_N19(clk_48Mhz__L6_N19), 
	.clk_48Mhz__L6_N2(clk_48Mhz__L6_N2), 
	.clk_48Mhz__L6_N20(clk_48Mhz__L6_N20), 
	.clk_48Mhz__L6_N21(clk_48Mhz__L6_N21), 
	.clk_48Mhz__L6_N22(clk_48Mhz__L6_N22), 
	.clk_48Mhz__L6_N23(clk_48Mhz__L6_N23), 
	.clk_48Mhz__L6_N24(clk_48Mhz__L6_N24), 
	.clk_48Mhz__L6_N25(clk_48Mhz__L6_N25), 
	.clk_48Mhz__L6_N26(clk_48Mhz__L6_N26), 
	.clk_48Mhz__L6_N27(clk_48Mhz__L6_N27), 
	.clk_48Mhz__L6_N28(clk_48Mhz__L6_N28), 
	.clk_48Mhz__L6_N29(clk_48Mhz__L6_N29), 
	.clk_48Mhz__L6_N3(clk_48Mhz__L6_N3), 
	.clk_48Mhz__L6_N30(clk_48Mhz__L6_N30), 
	.clk_48Mhz__L6_N31(clk_48Mhz__L6_N31), 
	.clk_48Mhz__L6_N32(clk_48Mhz__L6_N32), 
	.clk_48Mhz__L6_N33(clk_48Mhz__L6_N33), 
	.clk_48Mhz__L6_N34(clk_48Mhz__L6_N34), 
	.clk_48Mhz__L6_N35(clk_48Mhz__L6_N35), 
	.clk_48Mhz__L6_N36(clk_48Mhz__L6_N36), 
	.clk_48Mhz__L6_N37(clk_48Mhz__L6_N37), 
	.clk_48Mhz__L6_N38(clk_48Mhz__L6_N38), 
	.clk_48Mhz__L6_N39(clk_48Mhz__L6_N39), 
	.clk_48Mhz__L6_N4(clk_48Mhz__L6_N4), 
	.clk_48Mhz__L6_N40(clk_48Mhz__L6_N40), 
	.clk_48Mhz__L6_N41(clk_48Mhz__L6_N41), 
	.clk_48Mhz__L6_N42(clk_48Mhz__L6_N42), 
	.clk_48Mhz__L6_N43(clk_48Mhz__L6_N43), 
	.clk_48Mhz__L6_N44(clk_48Mhz__L6_N44), 
	.clk_48Mhz__L6_N45(clk_48Mhz__L6_N45), 
	.clk_48Mhz__L6_N46(clk_48Mhz__L6_N46), 
	.clk_48Mhz__L6_N47(clk_48Mhz__L6_N47), 
	.clk_48Mhz__L6_N5(clk_48Mhz__L6_N5), 
	.clk_48Mhz__L6_N6(clk_48Mhz__L6_N6), 
	.clk_48Mhz__L6_N7(clk_48Mhz__L6_N7), 
	.clk_48Mhz__L6_N8(clk_48Mhz__L6_N8), 
	.clk_48Mhz__L6_N9(clk_48Mhz__L6_N9));
   reg_in reg_in (.reset_n(FE_OFN37_reset_n), 
	.clk_48Mhz(clk_48Mhz__L6_N0), 
	.plain_byte_in(plain_byte_in), 
	.plain_byte_valid(plain_byte_valid), 
	.plain_finish(plain_finish), 
	.plain_key_out(Din), 
	.FE_OFN38_reset_n(FE_OFN38_reset_n), 
	.FE_OFN39_reset_n(FE_OFN39_reset_n), 
	.FE_OFN40_reset_n(FE_OFN40_reset_n), 
	.FE_OFN42_reset_n(FE_OFN42_reset_n), 
	.FE_OFN43_reset_n(FE_OFN43_reset_n), 
	.FE_OFN44_reset_n(FE_OFN44_reset_n), 
	.FE_OFN45_reset_n(FE_OFN45_reset_n), 
	.FE_OFN47_reset_n(FE_OFN47_reset_n), 
	.FE_OFN49_reset_n(FE_OFN49_reset_n), 
	.FE_OFN50_reset_n(FE_OFN50_reset_n), 
	.FE_OFN51_reset_n(FE_OFN51_reset_n), 
	.FE_OFN55_reset_n(FE_OFN55_reset_n), 
	.FE_OFN56_reset_n(FE_OFN56_reset_n), 
	.FE_OFN58_reset_n(FE_OFN58_reset_n), 
	.clk_48Mhz__L6_N1(clk_48Mhz__L6_N1), 
	.clk_48Mhz__L6_N10(clk_48Mhz__L6_N10), 
	.clk_48Mhz__L6_N11(clk_48Mhz__L6_N11), 
	.clk_48Mhz__L6_N14(clk_48Mhz__L6_N14), 
	.clk_48Mhz__L6_N15(clk_48Mhz__L6_N15), 
	.clk_48Mhz__L6_N2(clk_48Mhz__L6_N2), 
	.clk_48Mhz__L6_N20(clk_48Mhz__L6_N20), 
	.clk_48Mhz__L6_N21(clk_48Mhz__L6_N21), 
	.clk_48Mhz__L6_N23(clk_48Mhz__L6_N23), 
	.clk_48Mhz__L6_N25(clk_48Mhz__L6_N25), 
	.clk_48Mhz__L6_N27(clk_48Mhz__L6_N27), 
	.clk_48Mhz__L6_N28(clk_48Mhz__L6_N28), 
	.clk_48Mhz__L6_N29(clk_48Mhz__L6_N29), 
	.clk_48Mhz__L6_N35(clk_48Mhz__L6_N35), 
	.clk_48Mhz__L6_N37(clk_48Mhz__L6_N37), 
	.clk_48Mhz__L6_N39(clk_48Mhz__L6_N39), 
	.clk_48Mhz__L6_N4(clk_48Mhz__L6_N4), 
	.clk_48Mhz__L6_N40(clk_48Mhz__L6_N40), 
	.clk_48Mhz__L6_N41(clk_48Mhz__L6_N41), 
	.clk_48Mhz__L6_N5(clk_48Mhz__L6_N5), 
	.clk_48Mhz__L6_N6(clk_48Mhz__L6_N6), 
	.clk_48Mhz__L6_N8(clk_48Mhz__L6_N8), 
	.clk_48Mhz__L6_N9(clk_48Mhz__L6_N9));
   reg_out reg_out (.clk_48Mhz(clk_48Mhz__L6_N38), 
	.reset_n(FE_OFN38_reset_n), 
	.ready(ready), 
	.empty(empty), 
	.cipher_text(Dout), 
	.cipher_byte(cipher_byte_out), 
	.cipher_byte_valid(cipher_byte_valid), 
	.FE_OFN39_reset_n(FE_OFN39_reset_n), 
	.FE_OFN46_reset_n(FE_OFN46_reset_n), 
	.FE_OFN50_reset_n(FE_OFN50_reset_n), 
	.FE_OFN53_reset_n(FE_OFN53_reset_n), 
	.FE_OFN54_reset_n(FE_OFN54_reset_n), 
	.FE_OFN55_reset_n(FE_OFN55_reset_n), 
	.clk_48Mhz__L6_N39(clk_48Mhz__L6_N39), 
	.clk_48Mhz__L6_N41(clk_48Mhz__L6_N41), 
	.clk_48Mhz__L6_N43(clk_48Mhz__L6_N43), 
	.clk_48Mhz__L6_N44(clk_48Mhz__L6_N44), 
	.clk_48Mhz__L6_N45(clk_48Mhz__L6_N45), 
	.clk_48Mhz__L6_N46(clk_48Mhz__L6_N46), 
	.clk_48Mhz__L6_N47(clk_48Mhz__L6_N47));
endmodule

